module matmul (clk,
    rst,
    a,
    b,
    x);
 input clk;
 input rst;
 input [255:0] a;
 input [63:0] b;
 output [63:0] x;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire _22140_;
 wire _22141_;
 wire _22142_;
 wire _22143_;
 wire _22144_;
 wire _22145_;
 wire _22146_;
 wire _22147_;
 wire _22148_;
 wire _22149_;
 wire _22150_;
 wire _22151_;
 wire _22152_;
 wire _22153_;
 wire _22154_;
 wire _22155_;
 wire _22156_;
 wire _22157_;
 wire _22158_;
 wire _22159_;
 wire _22160_;
 wire _22161_;
 wire _22162_;
 wire _22163_;
 wire _22164_;
 wire _22165_;
 wire _22166_;
 wire _22167_;
 wire _22168_;
 wire _22169_;
 wire _22170_;
 wire _22171_;
 wire _22172_;
 wire _22173_;
 wire _22174_;
 wire _22175_;
 wire _22176_;
 wire _22177_;
 wire _22178_;
 wire _22179_;
 wire _22180_;
 wire _22181_;
 wire _22182_;
 wire _22183_;
 wire _22184_;
 wire _22185_;
 wire _22186_;
 wire _22187_;
 wire _22188_;
 wire _22189_;
 wire _22190_;
 wire _22191_;
 wire _22192_;
 wire _22193_;
 wire _22194_;
 wire _22195_;
 wire _22196_;
 wire _22197_;
 wire _22198_;
 wire _22199_;
 wire _22200_;
 wire _22201_;
 wire _22202_;
 wire _22203_;
 wire _22204_;
 wire _22205_;
 wire _22206_;
 wire _22207_;
 wire _22208_;
 wire _22209_;
 wire _22210_;
 wire _22211_;
 wire _22212_;
 wire _22213_;
 wire _22214_;
 wire _22215_;
 wire _22216_;
 wire _22217_;
 wire _22218_;
 wire _22219_;
 wire _22220_;
 wire _22221_;
 wire _22222_;
 wire _22223_;
 wire _22224_;
 wire _22225_;
 wire _22226_;
 wire _22227_;
 wire _22228_;
 wire _22229_;
 wire _22230_;
 wire _22231_;
 wire _22232_;
 wire _22233_;
 wire _22234_;
 wire _22235_;
 wire _22236_;
 wire _22237_;
 wire _22238_;
 wire _22239_;
 wire _22240_;
 wire _22241_;
 wire _22242_;
 wire _22243_;
 wire _22244_;
 wire _22245_;
 wire _22246_;
 wire _22247_;
 wire _22248_;
 wire _22249_;
 wire _22250_;
 wire _22251_;
 wire _22252_;
 wire _22253_;
 wire _22254_;
 wire _22255_;
 wire _22256_;
 wire _22257_;
 wire _22258_;
 wire _22259_;
 wire _22260_;
 wire _22261_;
 wire _22262_;
 wire _22263_;
 wire _22264_;
 wire _22265_;
 wire _22266_;
 wire _22267_;
 wire _22268_;
 wire _22269_;
 wire _22270_;
 wire _22271_;
 wire _22272_;
 wire _22273_;
 wire _22274_;
 wire _22275_;
 wire _22276_;
 wire _22277_;
 wire _22278_;
 wire _22279_;
 wire _22280_;
 wire _22281_;
 wire _22282_;
 wire _22283_;
 wire _22284_;
 wire _22285_;
 wire _22286_;
 wire _22287_;
 wire _22288_;
 wire _22289_;
 wire _22290_;
 wire _22291_;
 wire _22292_;
 wire _22293_;
 wire _22294_;
 wire _22295_;
 wire _22296_;
 wire _22297_;
 wire _22298_;
 wire _22299_;
 wire _22300_;
 wire _22301_;
 wire _22302_;
 wire _22303_;
 wire _22304_;
 wire _22305_;
 wire _22306_;
 wire _22307_;
 wire _22308_;
 wire _22309_;
 wire _22310_;
 wire _22311_;
 wire _22312_;
 wire _22313_;
 wire _22314_;
 wire _22315_;
 wire _22316_;
 wire _22317_;
 wire _22318_;
 wire _22319_;
 wire _22320_;
 wire _22321_;
 wire _22322_;
 wire _22323_;
 wire _22324_;
 wire _22325_;
 wire _22326_;
 wire _22327_;
 wire _22328_;
 wire _22329_;
 wire _22330_;
 wire _22331_;
 wire _22332_;
 wire _22333_;
 wire _22334_;
 wire _22335_;
 wire _22336_;
 wire _22337_;
 wire _22338_;
 wire _22339_;
 wire _22340_;
 wire _22341_;
 wire _22342_;
 wire _22343_;
 wire _22344_;
 wire _22345_;
 wire _22346_;
 wire _22347_;
 wire _22348_;
 wire _22349_;
 wire _22350_;
 wire _22351_;
 wire _22352_;
 wire _22353_;
 wire _22354_;
 wire _22355_;
 wire _22356_;
 wire _22357_;
 wire _22358_;
 wire _22359_;
 wire _22360_;
 wire _22361_;
 wire _22362_;
 wire _22363_;
 wire _22364_;
 wire _22365_;
 wire _22366_;
 wire _22367_;
 wire _22368_;
 wire _22369_;
 wire _22370_;
 wire _22371_;
 wire _22372_;
 wire _22373_;
 wire _22374_;
 wire _22375_;
 wire _22376_;
 wire _22377_;
 wire _22378_;
 wire _22379_;
 wire _22380_;
 wire _22381_;
 wire _22382_;
 wire _22383_;
 wire _22384_;
 wire _22385_;
 wire _22386_;
 wire _22387_;
 wire _22388_;
 wire _22389_;
 wire _22390_;
 wire _22391_;
 wire _22392_;
 wire _22393_;
 wire _22394_;
 wire _22395_;
 wire _22396_;
 wire _22397_;
 wire _22398_;
 wire _22399_;
 wire _22400_;
 wire _22401_;
 wire _22402_;
 wire _22403_;
 wire _22404_;
 wire _22405_;
 wire _22406_;
 wire _22407_;
 wire _22408_;
 wire _22409_;
 wire _22410_;
 wire _22411_;
 wire _22412_;
 wire _22413_;
 wire _22414_;
 wire _22415_;
 wire _22416_;
 wire _22417_;
 wire _22418_;
 wire _22419_;
 wire _22420_;
 wire _22421_;
 wire _22422_;
 wire _22423_;
 wire _22424_;
 wire _22425_;
 wire _22426_;
 wire _22427_;
 wire _22428_;
 wire _22429_;
 wire _22430_;
 wire _22431_;
 wire _22432_;
 wire _22433_;
 wire _22434_;
 wire _22435_;
 wire _22436_;
 wire _22437_;
 wire _22438_;
 wire _22439_;
 wire _22440_;
 wire _22441_;
 wire _22442_;
 wire _22443_;
 wire _22444_;
 wire _22445_;
 wire _22446_;
 wire _22447_;
 wire _22448_;
 wire _22449_;
 wire _22450_;
 wire _22451_;
 wire _22452_;
 wire _22453_;
 wire _22454_;
 wire _22455_;
 wire _22456_;
 wire _22457_;
 wire _22458_;
 wire _22459_;
 wire _22460_;
 wire _22461_;
 wire _22462_;
 wire _22463_;
 wire _22464_;
 wire _22465_;
 wire _22466_;
 wire _22467_;
 wire _22468_;
 wire _22469_;
 wire _22470_;
 wire _22471_;
 wire _22472_;
 wire _22473_;
 wire _22474_;
 wire _22475_;
 wire _22476_;
 wire _22477_;
 wire _22478_;
 wire _22479_;
 wire _22480_;
 wire _22481_;
 wire _22482_;
 wire _22483_;
 wire _22484_;
 wire _22485_;
 wire _22486_;
 wire _22487_;
 wire _22488_;
 wire _22489_;
 wire _22490_;
 wire _22491_;
 wire _22492_;
 wire _22493_;
 wire _22494_;
 wire _22495_;
 wire _22496_;
 wire _22497_;
 wire _22498_;
 wire _22499_;
 wire _22500_;
 wire _22501_;
 wire _22502_;
 wire _22503_;
 wire _22504_;
 wire _22505_;
 wire _22506_;
 wire _22507_;
 wire _22508_;
 wire _22509_;
 wire _22510_;
 wire _22511_;
 wire _22512_;
 wire _22513_;
 wire _22514_;
 wire _22515_;
 wire _22516_;
 wire _22517_;
 wire _22518_;
 wire _22519_;
 wire _22520_;
 wire _22521_;
 wire _22522_;
 wire _22523_;
 wire _22524_;
 wire _22525_;
 wire _22526_;
 wire _22527_;
 wire _22528_;
 wire _22529_;
 wire _22530_;
 wire _22531_;
 wire _22532_;
 wire _22533_;
 wire _22534_;
 wire _22535_;
 wire _22536_;
 wire _22537_;
 wire _22538_;
 wire _22539_;
 wire _22540_;
 wire _22541_;
 wire _22542_;
 wire _22543_;
 wire _22544_;
 wire _22545_;
 wire _22546_;
 wire _22547_;
 wire _22548_;
 wire _22549_;
 wire _22550_;
 wire _22551_;
 wire _22552_;
 wire _22553_;
 wire _22554_;
 wire _22555_;
 wire _22556_;
 wire _22557_;
 wire _22558_;
 wire clknet_leaf_0_clk;
 wire \g_reduce0[0].adder.a[0] ;
 wire \g_reduce0[0].adder.a[10] ;
 wire \g_reduce0[0].adder.a[11] ;
 wire \g_reduce0[0].adder.a[12] ;
 wire \g_reduce0[0].adder.a[13] ;
 wire \g_reduce0[0].adder.a[14] ;
 wire \g_reduce0[0].adder.a[15] ;
 wire \g_reduce0[0].adder.a[1] ;
 wire \g_reduce0[0].adder.a[2] ;
 wire \g_reduce0[0].adder.a[3] ;
 wire \g_reduce0[0].adder.a[4] ;
 wire \g_reduce0[0].adder.a[5] ;
 wire \g_reduce0[0].adder.a[6] ;
 wire \g_reduce0[0].adder.a[7] ;
 wire \g_reduce0[0].adder.a[8] ;
 wire \g_reduce0[0].adder.a[9] ;
 wire \g_reduce0[0].adder.b[0] ;
 wire \g_reduce0[0].adder.b[10] ;
 wire \g_reduce0[0].adder.b[11] ;
 wire \g_reduce0[0].adder.b[12] ;
 wire \g_reduce0[0].adder.b[13] ;
 wire \g_reduce0[0].adder.b[14] ;
 wire \g_reduce0[0].adder.b[15] ;
 wire \g_reduce0[0].adder.b[1] ;
 wire \g_reduce0[0].adder.b[2] ;
 wire \g_reduce0[0].adder.b[3] ;
 wire \g_reduce0[0].adder.b[4] ;
 wire \g_reduce0[0].adder.b[5] ;
 wire \g_reduce0[0].adder.b[6] ;
 wire \g_reduce0[0].adder.b[7] ;
 wire \g_reduce0[0].adder.b[8] ;
 wire \g_reduce0[0].adder.b[9] ;
 wire \g_reduce0[0].adder.x[0] ;
 wire \g_reduce0[0].adder.x[10] ;
 wire \g_reduce0[0].adder.x[11] ;
 wire \g_reduce0[0].adder.x[12] ;
 wire \g_reduce0[0].adder.x[13] ;
 wire \g_reduce0[0].adder.x[14] ;
 wire \g_reduce0[0].adder.x[15] ;
 wire \g_reduce0[0].adder.x[1] ;
 wire \g_reduce0[0].adder.x[2] ;
 wire \g_reduce0[0].adder.x[3] ;
 wire \g_reduce0[0].adder.x[4] ;
 wire \g_reduce0[0].adder.x[5] ;
 wire \g_reduce0[0].adder.x[6] ;
 wire \g_reduce0[0].adder.x[7] ;
 wire \g_reduce0[0].adder.x[8] ;
 wire \g_reduce0[0].adder.x[9] ;
 wire \g_reduce0[10].adder.a[0] ;
 wire \g_reduce0[10].adder.a[10] ;
 wire \g_reduce0[10].adder.a[11] ;
 wire \g_reduce0[10].adder.a[12] ;
 wire \g_reduce0[10].adder.a[13] ;
 wire \g_reduce0[10].adder.a[14] ;
 wire \g_reduce0[10].adder.a[15] ;
 wire \g_reduce0[10].adder.a[1] ;
 wire \g_reduce0[10].adder.a[2] ;
 wire \g_reduce0[10].adder.a[3] ;
 wire \g_reduce0[10].adder.a[4] ;
 wire \g_reduce0[10].adder.a[5] ;
 wire \g_reduce0[10].adder.a[6] ;
 wire \g_reduce0[10].adder.a[7] ;
 wire \g_reduce0[10].adder.a[8] ;
 wire \g_reduce0[10].adder.a[9] ;
 wire \g_reduce0[10].adder.b[0] ;
 wire \g_reduce0[10].adder.b[10] ;
 wire \g_reduce0[10].adder.b[11] ;
 wire \g_reduce0[10].adder.b[12] ;
 wire \g_reduce0[10].adder.b[13] ;
 wire \g_reduce0[10].adder.b[14] ;
 wire \g_reduce0[10].adder.b[15] ;
 wire \g_reduce0[10].adder.b[1] ;
 wire \g_reduce0[10].adder.b[2] ;
 wire \g_reduce0[10].adder.b[3] ;
 wire \g_reduce0[10].adder.b[4] ;
 wire \g_reduce0[10].adder.b[5] ;
 wire \g_reduce0[10].adder.b[6] ;
 wire \g_reduce0[10].adder.b[7] ;
 wire \g_reduce0[10].adder.b[8] ;
 wire \g_reduce0[10].adder.b[9] ;
 wire \g_reduce0[10].adder.x[0] ;
 wire \g_reduce0[10].adder.x[10] ;
 wire \g_reduce0[10].adder.x[11] ;
 wire \g_reduce0[10].adder.x[12] ;
 wire \g_reduce0[10].adder.x[13] ;
 wire \g_reduce0[10].adder.x[14] ;
 wire \g_reduce0[10].adder.x[15] ;
 wire \g_reduce0[10].adder.x[1] ;
 wire \g_reduce0[10].adder.x[2] ;
 wire \g_reduce0[10].adder.x[3] ;
 wire \g_reduce0[10].adder.x[4] ;
 wire \g_reduce0[10].adder.x[5] ;
 wire \g_reduce0[10].adder.x[6] ;
 wire \g_reduce0[10].adder.x[7] ;
 wire \g_reduce0[10].adder.x[8] ;
 wire \g_reduce0[10].adder.x[9] ;
 wire \g_reduce0[12].adder.a[0] ;
 wire \g_reduce0[12].adder.a[10] ;
 wire \g_reduce0[12].adder.a[11] ;
 wire \g_reduce0[12].adder.a[12] ;
 wire \g_reduce0[12].adder.a[13] ;
 wire \g_reduce0[12].adder.a[14] ;
 wire \g_reduce0[12].adder.a[15] ;
 wire \g_reduce0[12].adder.a[1] ;
 wire \g_reduce0[12].adder.a[2] ;
 wire \g_reduce0[12].adder.a[3] ;
 wire \g_reduce0[12].adder.a[4] ;
 wire \g_reduce0[12].adder.a[5] ;
 wire \g_reduce0[12].adder.a[6] ;
 wire \g_reduce0[12].adder.a[7] ;
 wire \g_reduce0[12].adder.a[8] ;
 wire \g_reduce0[12].adder.a[9] ;
 wire \g_reduce0[12].adder.b[0] ;
 wire \g_reduce0[12].adder.b[10] ;
 wire \g_reduce0[12].adder.b[11] ;
 wire \g_reduce0[12].adder.b[12] ;
 wire \g_reduce0[12].adder.b[13] ;
 wire \g_reduce0[12].adder.b[14] ;
 wire \g_reduce0[12].adder.b[15] ;
 wire \g_reduce0[12].adder.b[1] ;
 wire \g_reduce0[12].adder.b[2] ;
 wire \g_reduce0[12].adder.b[3] ;
 wire \g_reduce0[12].adder.b[4] ;
 wire \g_reduce0[12].adder.b[5] ;
 wire \g_reduce0[12].adder.b[6] ;
 wire \g_reduce0[12].adder.b[7] ;
 wire \g_reduce0[12].adder.b[8] ;
 wire \g_reduce0[12].adder.b[9] ;
 wire \g_reduce0[12].adder.x[0] ;
 wire \g_reduce0[12].adder.x[10] ;
 wire \g_reduce0[12].adder.x[11] ;
 wire \g_reduce0[12].adder.x[12] ;
 wire \g_reduce0[12].adder.x[13] ;
 wire \g_reduce0[12].adder.x[14] ;
 wire \g_reduce0[12].adder.x[15] ;
 wire \g_reduce0[12].adder.x[1] ;
 wire \g_reduce0[12].adder.x[2] ;
 wire \g_reduce0[12].adder.x[3] ;
 wire \g_reduce0[12].adder.x[4] ;
 wire \g_reduce0[12].adder.x[5] ;
 wire \g_reduce0[12].adder.x[6] ;
 wire \g_reduce0[12].adder.x[7] ;
 wire \g_reduce0[12].adder.x[8] ;
 wire \g_reduce0[12].adder.x[9] ;
 wire \g_reduce0[14].adder.a[0] ;
 wire \g_reduce0[14].adder.a[10] ;
 wire \g_reduce0[14].adder.a[11] ;
 wire \g_reduce0[14].adder.a[12] ;
 wire \g_reduce0[14].adder.a[13] ;
 wire \g_reduce0[14].adder.a[14] ;
 wire \g_reduce0[14].adder.a[15] ;
 wire \g_reduce0[14].adder.a[1] ;
 wire \g_reduce0[14].adder.a[2] ;
 wire \g_reduce0[14].adder.a[3] ;
 wire \g_reduce0[14].adder.a[4] ;
 wire \g_reduce0[14].adder.a[5] ;
 wire \g_reduce0[14].adder.a[6] ;
 wire \g_reduce0[14].adder.a[7] ;
 wire \g_reduce0[14].adder.a[8] ;
 wire \g_reduce0[14].adder.a[9] ;
 wire \g_reduce0[14].adder.b[0] ;
 wire \g_reduce0[14].adder.b[10] ;
 wire \g_reduce0[14].adder.b[11] ;
 wire \g_reduce0[14].adder.b[12] ;
 wire \g_reduce0[14].adder.b[13] ;
 wire \g_reduce0[14].adder.b[14] ;
 wire \g_reduce0[14].adder.b[15] ;
 wire \g_reduce0[14].adder.b[1] ;
 wire \g_reduce0[14].adder.b[2] ;
 wire \g_reduce0[14].adder.b[3] ;
 wire \g_reduce0[14].adder.b[4] ;
 wire \g_reduce0[14].adder.b[5] ;
 wire \g_reduce0[14].adder.b[6] ;
 wire \g_reduce0[14].adder.b[7] ;
 wire \g_reduce0[14].adder.b[8] ;
 wire \g_reduce0[14].adder.b[9] ;
 wire \g_reduce0[14].adder.x[0] ;
 wire \g_reduce0[14].adder.x[10] ;
 wire \g_reduce0[14].adder.x[11] ;
 wire \g_reduce0[14].adder.x[12] ;
 wire \g_reduce0[14].adder.x[13] ;
 wire \g_reduce0[14].adder.x[14] ;
 wire \g_reduce0[14].adder.x[15] ;
 wire \g_reduce0[14].adder.x[1] ;
 wire \g_reduce0[14].adder.x[2] ;
 wire \g_reduce0[14].adder.x[3] ;
 wire \g_reduce0[14].adder.x[4] ;
 wire \g_reduce0[14].adder.x[5] ;
 wire \g_reduce0[14].adder.x[6] ;
 wire \g_reduce0[14].adder.x[7] ;
 wire \g_reduce0[14].adder.x[8] ;
 wire \g_reduce0[14].adder.x[9] ;
 wire \g_reduce0[2].adder.a[0] ;
 wire \g_reduce0[2].adder.a[10] ;
 wire \g_reduce0[2].adder.a[11] ;
 wire \g_reduce0[2].adder.a[12] ;
 wire \g_reduce0[2].adder.a[13] ;
 wire \g_reduce0[2].adder.a[14] ;
 wire \g_reduce0[2].adder.a[15] ;
 wire \g_reduce0[2].adder.a[1] ;
 wire \g_reduce0[2].adder.a[2] ;
 wire \g_reduce0[2].adder.a[3] ;
 wire \g_reduce0[2].adder.a[4] ;
 wire \g_reduce0[2].adder.a[5] ;
 wire \g_reduce0[2].adder.a[6] ;
 wire \g_reduce0[2].adder.a[7] ;
 wire \g_reduce0[2].adder.a[8] ;
 wire \g_reduce0[2].adder.a[9] ;
 wire \g_reduce0[2].adder.b[0] ;
 wire \g_reduce0[2].adder.b[10] ;
 wire \g_reduce0[2].adder.b[11] ;
 wire \g_reduce0[2].adder.b[12] ;
 wire \g_reduce0[2].adder.b[13] ;
 wire \g_reduce0[2].adder.b[14] ;
 wire \g_reduce0[2].adder.b[15] ;
 wire \g_reduce0[2].adder.b[1] ;
 wire \g_reduce0[2].adder.b[2] ;
 wire \g_reduce0[2].adder.b[3] ;
 wire \g_reduce0[2].adder.b[4] ;
 wire \g_reduce0[2].adder.b[5] ;
 wire \g_reduce0[2].adder.b[6] ;
 wire \g_reduce0[2].adder.b[7] ;
 wire \g_reduce0[2].adder.b[8] ;
 wire \g_reduce0[2].adder.b[9] ;
 wire \g_reduce0[2].adder.x[0] ;
 wire \g_reduce0[2].adder.x[10] ;
 wire \g_reduce0[2].adder.x[11] ;
 wire \g_reduce0[2].adder.x[12] ;
 wire \g_reduce0[2].adder.x[13] ;
 wire \g_reduce0[2].adder.x[14] ;
 wire \g_reduce0[2].adder.x[15] ;
 wire \g_reduce0[2].adder.x[1] ;
 wire \g_reduce0[2].adder.x[2] ;
 wire \g_reduce0[2].adder.x[3] ;
 wire \g_reduce0[2].adder.x[4] ;
 wire \g_reduce0[2].adder.x[5] ;
 wire \g_reduce0[2].adder.x[6] ;
 wire \g_reduce0[2].adder.x[7] ;
 wire \g_reduce0[2].adder.x[8] ;
 wire \g_reduce0[2].adder.x[9] ;
 wire \g_reduce0[4].adder.a[0] ;
 wire \g_reduce0[4].adder.a[10] ;
 wire \g_reduce0[4].adder.a[11] ;
 wire \g_reduce0[4].adder.a[12] ;
 wire \g_reduce0[4].adder.a[13] ;
 wire \g_reduce0[4].adder.a[14] ;
 wire \g_reduce0[4].adder.a[15] ;
 wire \g_reduce0[4].adder.a[1] ;
 wire \g_reduce0[4].adder.a[2] ;
 wire \g_reduce0[4].adder.a[3] ;
 wire \g_reduce0[4].adder.a[4] ;
 wire \g_reduce0[4].adder.a[5] ;
 wire \g_reduce0[4].adder.a[6] ;
 wire \g_reduce0[4].adder.a[7] ;
 wire \g_reduce0[4].adder.a[8] ;
 wire \g_reduce0[4].adder.a[9] ;
 wire \g_reduce0[4].adder.b[0] ;
 wire \g_reduce0[4].adder.b[10] ;
 wire \g_reduce0[4].adder.b[11] ;
 wire \g_reduce0[4].adder.b[12] ;
 wire \g_reduce0[4].adder.b[13] ;
 wire \g_reduce0[4].adder.b[14] ;
 wire \g_reduce0[4].adder.b[15] ;
 wire \g_reduce0[4].adder.b[1] ;
 wire \g_reduce0[4].adder.b[2] ;
 wire \g_reduce0[4].adder.b[3] ;
 wire \g_reduce0[4].adder.b[4] ;
 wire \g_reduce0[4].adder.b[5] ;
 wire \g_reduce0[4].adder.b[6] ;
 wire \g_reduce0[4].adder.b[7] ;
 wire \g_reduce0[4].adder.b[8] ;
 wire \g_reduce0[4].adder.b[9] ;
 wire \g_reduce0[4].adder.x[0] ;
 wire \g_reduce0[4].adder.x[10] ;
 wire \g_reduce0[4].adder.x[11] ;
 wire \g_reduce0[4].adder.x[12] ;
 wire \g_reduce0[4].adder.x[13] ;
 wire \g_reduce0[4].adder.x[14] ;
 wire \g_reduce0[4].adder.x[15] ;
 wire \g_reduce0[4].adder.x[1] ;
 wire \g_reduce0[4].adder.x[2] ;
 wire \g_reduce0[4].adder.x[3] ;
 wire \g_reduce0[4].adder.x[4] ;
 wire \g_reduce0[4].adder.x[5] ;
 wire \g_reduce0[4].adder.x[6] ;
 wire \g_reduce0[4].adder.x[7] ;
 wire \g_reduce0[4].adder.x[8] ;
 wire \g_reduce0[4].adder.x[9] ;
 wire \g_reduce0[6].adder.a[0] ;
 wire \g_reduce0[6].adder.a[10] ;
 wire \g_reduce0[6].adder.a[11] ;
 wire \g_reduce0[6].adder.a[12] ;
 wire \g_reduce0[6].adder.a[13] ;
 wire \g_reduce0[6].adder.a[14] ;
 wire \g_reduce0[6].adder.a[15] ;
 wire \g_reduce0[6].adder.a[1] ;
 wire \g_reduce0[6].adder.a[2] ;
 wire \g_reduce0[6].adder.a[3] ;
 wire \g_reduce0[6].adder.a[4] ;
 wire \g_reduce0[6].adder.a[5] ;
 wire \g_reduce0[6].adder.a[6] ;
 wire \g_reduce0[6].adder.a[7] ;
 wire \g_reduce0[6].adder.a[8] ;
 wire \g_reduce0[6].adder.a[9] ;
 wire \g_reduce0[6].adder.b[0] ;
 wire \g_reduce0[6].adder.b[10] ;
 wire \g_reduce0[6].adder.b[11] ;
 wire \g_reduce0[6].adder.b[12] ;
 wire \g_reduce0[6].adder.b[13] ;
 wire \g_reduce0[6].adder.b[14] ;
 wire \g_reduce0[6].adder.b[15] ;
 wire \g_reduce0[6].adder.b[1] ;
 wire \g_reduce0[6].adder.b[2] ;
 wire \g_reduce0[6].adder.b[3] ;
 wire \g_reduce0[6].adder.b[4] ;
 wire \g_reduce0[6].adder.b[5] ;
 wire \g_reduce0[6].adder.b[6] ;
 wire \g_reduce0[6].adder.b[7] ;
 wire \g_reduce0[6].adder.b[8] ;
 wire \g_reduce0[6].adder.b[9] ;
 wire \g_reduce0[6].adder.x[0] ;
 wire \g_reduce0[6].adder.x[10] ;
 wire \g_reduce0[6].adder.x[11] ;
 wire \g_reduce0[6].adder.x[12] ;
 wire \g_reduce0[6].adder.x[13] ;
 wire \g_reduce0[6].adder.x[14] ;
 wire \g_reduce0[6].adder.x[15] ;
 wire \g_reduce0[6].adder.x[1] ;
 wire \g_reduce0[6].adder.x[2] ;
 wire \g_reduce0[6].adder.x[3] ;
 wire \g_reduce0[6].adder.x[4] ;
 wire \g_reduce0[6].adder.x[5] ;
 wire \g_reduce0[6].adder.x[6] ;
 wire \g_reduce0[6].adder.x[7] ;
 wire \g_reduce0[6].adder.x[8] ;
 wire \g_reduce0[6].adder.x[9] ;
 wire \g_reduce0[8].adder.a[0] ;
 wire \g_reduce0[8].adder.a[10] ;
 wire \g_reduce0[8].adder.a[11] ;
 wire \g_reduce0[8].adder.a[12] ;
 wire \g_reduce0[8].adder.a[13] ;
 wire \g_reduce0[8].adder.a[14] ;
 wire \g_reduce0[8].adder.a[15] ;
 wire \g_reduce0[8].adder.a[1] ;
 wire \g_reduce0[8].adder.a[2] ;
 wire \g_reduce0[8].adder.a[3] ;
 wire \g_reduce0[8].adder.a[4] ;
 wire \g_reduce0[8].adder.a[5] ;
 wire \g_reduce0[8].adder.a[6] ;
 wire \g_reduce0[8].adder.a[7] ;
 wire \g_reduce0[8].adder.a[8] ;
 wire \g_reduce0[8].adder.a[9] ;
 wire \g_reduce0[8].adder.b[0] ;
 wire \g_reduce0[8].adder.b[10] ;
 wire \g_reduce0[8].adder.b[11] ;
 wire \g_reduce0[8].adder.b[12] ;
 wire \g_reduce0[8].adder.b[13] ;
 wire \g_reduce0[8].adder.b[14] ;
 wire \g_reduce0[8].adder.b[15] ;
 wire \g_reduce0[8].adder.b[1] ;
 wire \g_reduce0[8].adder.b[2] ;
 wire \g_reduce0[8].adder.b[3] ;
 wire \g_reduce0[8].adder.b[4] ;
 wire \g_reduce0[8].adder.b[5] ;
 wire \g_reduce0[8].adder.b[6] ;
 wire \g_reduce0[8].adder.b[7] ;
 wire \g_reduce0[8].adder.b[8] ;
 wire \g_reduce0[8].adder.b[9] ;
 wire \g_reduce0[8].adder.x[0] ;
 wire \g_reduce0[8].adder.x[10] ;
 wire \g_reduce0[8].adder.x[11] ;
 wire \g_reduce0[8].adder.x[12] ;
 wire \g_reduce0[8].adder.x[13] ;
 wire \g_reduce0[8].adder.x[14] ;
 wire \g_reduce0[8].adder.x[15] ;
 wire \g_reduce0[8].adder.x[1] ;
 wire \g_reduce0[8].adder.x[2] ;
 wire \g_reduce0[8].adder.x[3] ;
 wire \g_reduce0[8].adder.x[4] ;
 wire \g_reduce0[8].adder.x[5] ;
 wire \g_reduce0[8].adder.x[6] ;
 wire \g_reduce0[8].adder.x[7] ;
 wire \g_reduce0[8].adder.x[8] ;
 wire \g_reduce0[8].adder.x[9] ;
 wire \g_row[0].g_col[0].mult.adder.a[0] ;
 wire \g_row[0].g_col[0].mult.adder.a[10] ;
 wire \g_row[0].g_col[0].mult.adder.a[11] ;
 wire \g_row[0].g_col[0].mult.adder.a[12] ;
 wire \g_row[0].g_col[0].mult.adder.a[13] ;
 wire \g_row[0].g_col[0].mult.adder.a[14] ;
 wire \g_row[0].g_col[0].mult.adder.a[15] ;
 wire \g_row[0].g_col[0].mult.adder.a[16] ;
 wire \g_row[0].g_col[0].mult.adder.a[17] ;
 wire \g_row[0].g_col[0].mult.adder.a[18] ;
 wire \g_row[0].g_col[0].mult.adder.a[19] ;
 wire \g_row[0].g_col[0].mult.adder.a[1] ;
 wire \g_row[0].g_col[0].mult.adder.a[20] ;
 wire \g_row[0].g_col[0].mult.adder.a[2] ;
 wire \g_row[0].g_col[0].mult.adder.a[3] ;
 wire \g_row[0].g_col[0].mult.adder.a[4] ;
 wire \g_row[0].g_col[0].mult.adder.a[5] ;
 wire \g_row[0].g_col[0].mult.adder.a[6] ;
 wire \g_row[0].g_col[0].mult.adder.a[7] ;
 wire \g_row[0].g_col[0].mult.adder.a[8] ;
 wire \g_row[0].g_col[0].mult.adder.a[9] ;
 wire \g_row[0].g_col[0].mult.adder.b[10] ;
 wire \g_row[0].g_col[0].mult.adder.b[11] ;
 wire \g_row[0].g_col[0].mult.adder.b[12] ;
 wire \g_row[0].g_col[0].mult.adder.b[13] ;
 wire \g_row[0].g_col[0].mult.adder.b[14] ;
 wire \g_row[0].g_col[0].mult.adder.b[15] ;
 wire \g_row[0].g_col[0].mult.adder.b[16] ;
 wire \g_row[0].g_col[0].mult.adder.b[17] ;
 wire \g_row[0].g_col[0].mult.adder.b[18] ;
 wire \g_row[0].g_col[0].mult.adder.b[19] ;
 wire \g_row[0].g_col[0].mult.adder.b[1] ;
 wire \g_row[0].g_col[0].mult.adder.b[20] ;
 wire \g_row[0].g_col[0].mult.adder.b[2] ;
 wire \g_row[0].g_col[0].mult.adder.b[3] ;
 wire \g_row[0].g_col[0].mult.adder.b[4] ;
 wire \g_row[0].g_col[0].mult.adder.b[5] ;
 wire \g_row[0].g_col[0].mult.adder.b[6] ;
 wire \g_row[0].g_col[0].mult.adder.b[7] ;
 wire \g_row[0].g_col[0].mult.adder.b[8] ;
 wire \g_row[0].g_col[0].mult.adder.b[9] ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.b ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.b ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.b ;
 wire \g_row[0].g_col[0].mult.sign ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[0] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[10] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[11] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[12] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[13] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[14] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[15] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[16] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[17] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[18] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[19] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[1] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[2] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[3] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[4] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[5] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[6] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[7] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[8] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t1[9] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[10] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[11] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[12] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[13] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[14] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[15] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[16] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[17] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[18] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[19] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[1] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[20] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[2] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[3] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[4] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[5] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[6] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[7] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[8] ;
 wire \g_row[0].g_col[0].mult.stage1.dadda.t2[9] ;
 wire \g_row[0].g_col[1].mult.adder.a[0] ;
 wire \g_row[0].g_col[1].mult.adder.a[10] ;
 wire \g_row[0].g_col[1].mult.adder.a[11] ;
 wire \g_row[0].g_col[1].mult.adder.a[12] ;
 wire \g_row[0].g_col[1].mult.adder.a[13] ;
 wire \g_row[0].g_col[1].mult.adder.a[14] ;
 wire \g_row[0].g_col[1].mult.adder.a[15] ;
 wire \g_row[0].g_col[1].mult.adder.a[16] ;
 wire \g_row[0].g_col[1].mult.adder.a[17] ;
 wire \g_row[0].g_col[1].mult.adder.a[18] ;
 wire \g_row[0].g_col[1].mult.adder.a[19] ;
 wire \g_row[0].g_col[1].mult.adder.a[1] ;
 wire \g_row[0].g_col[1].mult.adder.a[2] ;
 wire \g_row[0].g_col[1].mult.adder.a[3] ;
 wire \g_row[0].g_col[1].mult.adder.a[4] ;
 wire \g_row[0].g_col[1].mult.adder.a[5] ;
 wire \g_row[0].g_col[1].mult.adder.a[6] ;
 wire \g_row[0].g_col[1].mult.adder.a[7] ;
 wire \g_row[0].g_col[1].mult.adder.a[8] ;
 wire \g_row[0].g_col[1].mult.adder.a[9] ;
 wire \g_row[0].g_col[1].mult.adder.b[10] ;
 wire \g_row[0].g_col[1].mult.adder.b[11] ;
 wire \g_row[0].g_col[1].mult.adder.b[12] ;
 wire \g_row[0].g_col[1].mult.adder.b[13] ;
 wire \g_row[0].g_col[1].mult.adder.b[14] ;
 wire \g_row[0].g_col[1].mult.adder.b[15] ;
 wire \g_row[0].g_col[1].mult.adder.b[16] ;
 wire \g_row[0].g_col[1].mult.adder.b[17] ;
 wire \g_row[0].g_col[1].mult.adder.b[18] ;
 wire \g_row[0].g_col[1].mult.adder.b[19] ;
 wire \g_row[0].g_col[1].mult.adder.b[1] ;
 wire \g_row[0].g_col[1].mult.adder.b[20] ;
 wire \g_row[0].g_col[1].mult.adder.b[2] ;
 wire \g_row[0].g_col[1].mult.adder.b[3] ;
 wire \g_row[0].g_col[1].mult.adder.b[4] ;
 wire \g_row[0].g_col[1].mult.adder.b[5] ;
 wire \g_row[0].g_col[1].mult.adder.b[6] ;
 wire \g_row[0].g_col[1].mult.adder.b[7] ;
 wire \g_row[0].g_col[1].mult.adder.b[8] ;
 wire \g_row[0].g_col[1].mult.adder.b[9] ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.b ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.b ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.b ;
 wire \g_row[0].g_col[1].mult.sign ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[0] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[10] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[11] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[12] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[13] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[14] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[15] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[16] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[17] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[18] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[19] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[1] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[2] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[3] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[4] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[5] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[6] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[7] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[8] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t1[9] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[10] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[11] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[12] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[13] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[14] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[15] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[16] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[17] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[18] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[19] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[1] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[20] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[2] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[3] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[4] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[5] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[6] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[7] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[8] ;
 wire \g_row[0].g_col[1].mult.stage1.dadda.t2[9] ;
 wire \g_row[0].g_col[2].mult.adder.a[0] ;
 wire \g_row[0].g_col[2].mult.adder.a[10] ;
 wire \g_row[0].g_col[2].mult.adder.a[11] ;
 wire \g_row[0].g_col[2].mult.adder.a[12] ;
 wire \g_row[0].g_col[2].mult.adder.a[13] ;
 wire \g_row[0].g_col[2].mult.adder.a[14] ;
 wire \g_row[0].g_col[2].mult.adder.a[15] ;
 wire \g_row[0].g_col[2].mult.adder.a[16] ;
 wire \g_row[0].g_col[2].mult.adder.a[17] ;
 wire \g_row[0].g_col[2].mult.adder.a[18] ;
 wire \g_row[0].g_col[2].mult.adder.a[19] ;
 wire \g_row[0].g_col[2].mult.adder.a[1] ;
 wire \g_row[0].g_col[2].mult.adder.a[2] ;
 wire \g_row[0].g_col[2].mult.adder.a[3] ;
 wire \g_row[0].g_col[2].mult.adder.a[4] ;
 wire \g_row[0].g_col[2].mult.adder.a[5] ;
 wire \g_row[0].g_col[2].mult.adder.a[6] ;
 wire \g_row[0].g_col[2].mult.adder.a[7] ;
 wire \g_row[0].g_col[2].mult.adder.a[8] ;
 wire \g_row[0].g_col[2].mult.adder.a[9] ;
 wire \g_row[0].g_col[2].mult.adder.b[10] ;
 wire \g_row[0].g_col[2].mult.adder.b[11] ;
 wire \g_row[0].g_col[2].mult.adder.b[12] ;
 wire \g_row[0].g_col[2].mult.adder.b[13] ;
 wire \g_row[0].g_col[2].mult.adder.b[14] ;
 wire \g_row[0].g_col[2].mult.adder.b[15] ;
 wire \g_row[0].g_col[2].mult.adder.b[16] ;
 wire \g_row[0].g_col[2].mult.adder.b[17] ;
 wire \g_row[0].g_col[2].mult.adder.b[18] ;
 wire \g_row[0].g_col[2].mult.adder.b[19] ;
 wire \g_row[0].g_col[2].mult.adder.b[1] ;
 wire \g_row[0].g_col[2].mult.adder.b[20] ;
 wire \g_row[0].g_col[2].mult.adder.b[2] ;
 wire \g_row[0].g_col[2].mult.adder.b[3] ;
 wire \g_row[0].g_col[2].mult.adder.b[4] ;
 wire \g_row[0].g_col[2].mult.adder.b[5] ;
 wire \g_row[0].g_col[2].mult.adder.b[6] ;
 wire \g_row[0].g_col[2].mult.adder.b[7] ;
 wire \g_row[0].g_col[2].mult.adder.b[8] ;
 wire \g_row[0].g_col[2].mult.adder.b[9] ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.b ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.b ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.b ;
 wire \g_row[0].g_col[2].mult.sign ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[0] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[10] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[11] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[12] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[13] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[14] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[15] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[16] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[17] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[18] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[19] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[1] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[2] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[3] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[4] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[5] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[6] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[7] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[8] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t1[9] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[10] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[11] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[12] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[13] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[14] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[15] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[16] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[17] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[18] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[19] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[1] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[20] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[2] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[3] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[4] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[5] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[6] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[7] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[8] ;
 wire \g_row[0].g_col[2].mult.stage1.dadda.t2[9] ;
 wire \g_row[0].g_col[3].mult.adder.a[0] ;
 wire \g_row[0].g_col[3].mult.adder.a[10] ;
 wire \g_row[0].g_col[3].mult.adder.a[11] ;
 wire \g_row[0].g_col[3].mult.adder.a[12] ;
 wire \g_row[0].g_col[3].mult.adder.a[13] ;
 wire \g_row[0].g_col[3].mult.adder.a[14] ;
 wire \g_row[0].g_col[3].mult.adder.a[15] ;
 wire \g_row[0].g_col[3].mult.adder.a[16] ;
 wire \g_row[0].g_col[3].mult.adder.a[17] ;
 wire \g_row[0].g_col[3].mult.adder.a[18] ;
 wire \g_row[0].g_col[3].mult.adder.a[19] ;
 wire \g_row[0].g_col[3].mult.adder.a[1] ;
 wire \g_row[0].g_col[3].mult.adder.a[2] ;
 wire \g_row[0].g_col[3].mult.adder.a[3] ;
 wire \g_row[0].g_col[3].mult.adder.a[4] ;
 wire \g_row[0].g_col[3].mult.adder.a[5] ;
 wire \g_row[0].g_col[3].mult.adder.a[6] ;
 wire \g_row[0].g_col[3].mult.adder.a[7] ;
 wire \g_row[0].g_col[3].mult.adder.a[8] ;
 wire \g_row[0].g_col[3].mult.adder.a[9] ;
 wire \g_row[0].g_col[3].mult.adder.b[10] ;
 wire \g_row[0].g_col[3].mult.adder.b[11] ;
 wire \g_row[0].g_col[3].mult.adder.b[12] ;
 wire \g_row[0].g_col[3].mult.adder.b[13] ;
 wire \g_row[0].g_col[3].mult.adder.b[14] ;
 wire \g_row[0].g_col[3].mult.adder.b[15] ;
 wire \g_row[0].g_col[3].mult.adder.b[16] ;
 wire \g_row[0].g_col[3].mult.adder.b[17] ;
 wire \g_row[0].g_col[3].mult.adder.b[18] ;
 wire \g_row[0].g_col[3].mult.adder.b[19] ;
 wire \g_row[0].g_col[3].mult.adder.b[1] ;
 wire \g_row[0].g_col[3].mult.adder.b[20] ;
 wire \g_row[0].g_col[3].mult.adder.b[2] ;
 wire \g_row[0].g_col[3].mult.adder.b[3] ;
 wire \g_row[0].g_col[3].mult.adder.b[4] ;
 wire \g_row[0].g_col[3].mult.adder.b[5] ;
 wire \g_row[0].g_col[3].mult.adder.b[6] ;
 wire \g_row[0].g_col[3].mult.adder.b[7] ;
 wire \g_row[0].g_col[3].mult.adder.b[8] ;
 wire \g_row[0].g_col[3].mult.adder.b[9] ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.b ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.b ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.b ;
 wire \g_row[0].g_col[3].mult.sign ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[0] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[10] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[11] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[12] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[13] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[14] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[15] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[16] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[17] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[18] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[19] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[1] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[2] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[3] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[4] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[5] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[6] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[7] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[8] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t1[9] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[10] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[11] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[12] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[13] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[14] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[15] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[16] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[17] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[18] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[19] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[1] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[20] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[2] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[3] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[4] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[5] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[6] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[7] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[8] ;
 wire \g_row[0].g_col[3].mult.stage1.dadda.t2[9] ;
 wire \g_row[1].g_col[0].mult.adder.a[0] ;
 wire \g_row[1].g_col[0].mult.adder.a[10] ;
 wire \g_row[1].g_col[0].mult.adder.a[11] ;
 wire \g_row[1].g_col[0].mult.adder.a[12] ;
 wire \g_row[1].g_col[0].mult.adder.a[13] ;
 wire \g_row[1].g_col[0].mult.adder.a[14] ;
 wire \g_row[1].g_col[0].mult.adder.a[15] ;
 wire \g_row[1].g_col[0].mult.adder.a[16] ;
 wire \g_row[1].g_col[0].mult.adder.a[17] ;
 wire \g_row[1].g_col[0].mult.adder.a[18] ;
 wire \g_row[1].g_col[0].mult.adder.a[19] ;
 wire \g_row[1].g_col[0].mult.adder.a[1] ;
 wire \g_row[1].g_col[0].mult.adder.a[2] ;
 wire \g_row[1].g_col[0].mult.adder.a[3] ;
 wire \g_row[1].g_col[0].mult.adder.a[4] ;
 wire \g_row[1].g_col[0].mult.adder.a[5] ;
 wire \g_row[1].g_col[0].mult.adder.a[6] ;
 wire \g_row[1].g_col[0].mult.adder.a[7] ;
 wire \g_row[1].g_col[0].mult.adder.a[8] ;
 wire \g_row[1].g_col[0].mult.adder.a[9] ;
 wire \g_row[1].g_col[0].mult.adder.b[10] ;
 wire \g_row[1].g_col[0].mult.adder.b[11] ;
 wire \g_row[1].g_col[0].mult.adder.b[12] ;
 wire \g_row[1].g_col[0].mult.adder.b[13] ;
 wire \g_row[1].g_col[0].mult.adder.b[14] ;
 wire \g_row[1].g_col[0].mult.adder.b[15] ;
 wire \g_row[1].g_col[0].mult.adder.b[16] ;
 wire \g_row[1].g_col[0].mult.adder.b[17] ;
 wire \g_row[1].g_col[0].mult.adder.b[18] ;
 wire \g_row[1].g_col[0].mult.adder.b[19] ;
 wire \g_row[1].g_col[0].mult.adder.b[1] ;
 wire \g_row[1].g_col[0].mult.adder.b[20] ;
 wire \g_row[1].g_col[0].mult.adder.b[2] ;
 wire \g_row[1].g_col[0].mult.adder.b[3] ;
 wire \g_row[1].g_col[0].mult.adder.b[4] ;
 wire \g_row[1].g_col[0].mult.adder.b[5] ;
 wire \g_row[1].g_col[0].mult.adder.b[6] ;
 wire \g_row[1].g_col[0].mult.adder.b[7] ;
 wire \g_row[1].g_col[0].mult.adder.b[8] ;
 wire \g_row[1].g_col[0].mult.adder.b[9] ;
 wire \g_row[1].g_col[0].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[1].g_col[0].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[1].g_col[0].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[1].g_col[0].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[1].g_col[0].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[1].g_col[0].mult.sign ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[0] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[10] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[11] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[12] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[13] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[14] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[15] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[16] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[17] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[18] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[19] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[1] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[2] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[3] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[4] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[5] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[6] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[7] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[8] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t1[9] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[10] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[11] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[12] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[13] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[14] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[15] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[16] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[17] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[18] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[19] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[1] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[20] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[2] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[3] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[4] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[5] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[6] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[7] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[8] ;
 wire \g_row[1].g_col[0].mult.stage1.dadda.t2[9] ;
 wire \g_row[1].g_col[1].mult.adder.a[0] ;
 wire \g_row[1].g_col[1].mult.adder.a[10] ;
 wire \g_row[1].g_col[1].mult.adder.a[11] ;
 wire \g_row[1].g_col[1].mult.adder.a[12] ;
 wire \g_row[1].g_col[1].mult.adder.a[13] ;
 wire \g_row[1].g_col[1].mult.adder.a[14] ;
 wire \g_row[1].g_col[1].mult.adder.a[15] ;
 wire \g_row[1].g_col[1].mult.adder.a[16] ;
 wire \g_row[1].g_col[1].mult.adder.a[17] ;
 wire \g_row[1].g_col[1].mult.adder.a[18] ;
 wire \g_row[1].g_col[1].mult.adder.a[19] ;
 wire \g_row[1].g_col[1].mult.adder.a[1] ;
 wire \g_row[1].g_col[1].mult.adder.a[2] ;
 wire \g_row[1].g_col[1].mult.adder.a[3] ;
 wire \g_row[1].g_col[1].mult.adder.a[4] ;
 wire \g_row[1].g_col[1].mult.adder.a[5] ;
 wire \g_row[1].g_col[1].mult.adder.a[6] ;
 wire \g_row[1].g_col[1].mult.adder.a[7] ;
 wire \g_row[1].g_col[1].mult.adder.a[8] ;
 wire \g_row[1].g_col[1].mult.adder.a[9] ;
 wire \g_row[1].g_col[1].mult.adder.b[10] ;
 wire \g_row[1].g_col[1].mult.adder.b[11] ;
 wire \g_row[1].g_col[1].mult.adder.b[12] ;
 wire \g_row[1].g_col[1].mult.adder.b[13] ;
 wire \g_row[1].g_col[1].mult.adder.b[14] ;
 wire \g_row[1].g_col[1].mult.adder.b[15] ;
 wire \g_row[1].g_col[1].mult.adder.b[16] ;
 wire \g_row[1].g_col[1].mult.adder.b[17] ;
 wire \g_row[1].g_col[1].mult.adder.b[18] ;
 wire \g_row[1].g_col[1].mult.adder.b[19] ;
 wire \g_row[1].g_col[1].mult.adder.b[1] ;
 wire \g_row[1].g_col[1].mult.adder.b[20] ;
 wire \g_row[1].g_col[1].mult.adder.b[2] ;
 wire \g_row[1].g_col[1].mult.adder.b[3] ;
 wire \g_row[1].g_col[1].mult.adder.b[4] ;
 wire \g_row[1].g_col[1].mult.adder.b[5] ;
 wire \g_row[1].g_col[1].mult.adder.b[6] ;
 wire \g_row[1].g_col[1].mult.adder.b[7] ;
 wire \g_row[1].g_col[1].mult.adder.b[8] ;
 wire \g_row[1].g_col[1].mult.adder.b[9] ;
 wire \g_row[1].g_col[1].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[1].g_col[1].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[1].g_col[1].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[1].g_col[1].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[1].g_col[1].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[1].g_col[1].mult.sign ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[0] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[10] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[11] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[12] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[13] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[14] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[15] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[16] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[17] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[18] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[19] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[1] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[2] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[3] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[4] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[5] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[6] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[7] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[8] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t1[9] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[10] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[11] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[12] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[13] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[14] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[15] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[16] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[17] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[18] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[19] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[1] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[20] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[2] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[3] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[4] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[5] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[6] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[7] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[8] ;
 wire \g_row[1].g_col[1].mult.stage1.dadda.t2[9] ;
 wire \g_row[1].g_col[2].mult.adder.a[0] ;
 wire \g_row[1].g_col[2].mult.adder.a[10] ;
 wire \g_row[1].g_col[2].mult.adder.a[11] ;
 wire \g_row[1].g_col[2].mult.adder.a[12] ;
 wire \g_row[1].g_col[2].mult.adder.a[13] ;
 wire \g_row[1].g_col[2].mult.adder.a[14] ;
 wire \g_row[1].g_col[2].mult.adder.a[15] ;
 wire \g_row[1].g_col[2].mult.adder.a[16] ;
 wire \g_row[1].g_col[2].mult.adder.a[17] ;
 wire \g_row[1].g_col[2].mult.adder.a[18] ;
 wire \g_row[1].g_col[2].mult.adder.a[19] ;
 wire \g_row[1].g_col[2].mult.adder.a[1] ;
 wire \g_row[1].g_col[2].mult.adder.a[2] ;
 wire \g_row[1].g_col[2].mult.adder.a[3] ;
 wire \g_row[1].g_col[2].mult.adder.a[4] ;
 wire \g_row[1].g_col[2].mult.adder.a[5] ;
 wire \g_row[1].g_col[2].mult.adder.a[6] ;
 wire \g_row[1].g_col[2].mult.adder.a[7] ;
 wire \g_row[1].g_col[2].mult.adder.a[8] ;
 wire \g_row[1].g_col[2].mult.adder.a[9] ;
 wire \g_row[1].g_col[2].mult.adder.b[10] ;
 wire \g_row[1].g_col[2].mult.adder.b[11] ;
 wire \g_row[1].g_col[2].mult.adder.b[12] ;
 wire \g_row[1].g_col[2].mult.adder.b[13] ;
 wire \g_row[1].g_col[2].mult.adder.b[14] ;
 wire \g_row[1].g_col[2].mult.adder.b[15] ;
 wire \g_row[1].g_col[2].mult.adder.b[16] ;
 wire \g_row[1].g_col[2].mult.adder.b[17] ;
 wire \g_row[1].g_col[2].mult.adder.b[18] ;
 wire \g_row[1].g_col[2].mult.adder.b[19] ;
 wire \g_row[1].g_col[2].mult.adder.b[1] ;
 wire \g_row[1].g_col[2].mult.adder.b[20] ;
 wire \g_row[1].g_col[2].mult.adder.b[2] ;
 wire \g_row[1].g_col[2].mult.adder.b[3] ;
 wire \g_row[1].g_col[2].mult.adder.b[4] ;
 wire \g_row[1].g_col[2].mult.adder.b[5] ;
 wire \g_row[1].g_col[2].mult.adder.b[6] ;
 wire \g_row[1].g_col[2].mult.adder.b[7] ;
 wire \g_row[1].g_col[2].mult.adder.b[8] ;
 wire \g_row[1].g_col[2].mult.adder.b[9] ;
 wire \g_row[1].g_col[2].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[1].g_col[2].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[1].g_col[2].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[1].g_col[2].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[1].g_col[2].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[1].g_col[2].mult.sign ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[0] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[10] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[11] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[12] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[13] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[14] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[15] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[16] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[17] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[18] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[19] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[1] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[2] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[3] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[4] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[5] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[6] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[7] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[8] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t1[9] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[10] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[11] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[12] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[13] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[14] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[15] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[16] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[17] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[18] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[19] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[1] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[20] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[2] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[3] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[4] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[5] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[6] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[7] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[8] ;
 wire \g_row[1].g_col[2].mult.stage1.dadda.t2[9] ;
 wire \g_row[1].g_col[3].mult.adder.a[0] ;
 wire \g_row[1].g_col[3].mult.adder.a[10] ;
 wire \g_row[1].g_col[3].mult.adder.a[11] ;
 wire \g_row[1].g_col[3].mult.adder.a[12] ;
 wire \g_row[1].g_col[3].mult.adder.a[13] ;
 wire \g_row[1].g_col[3].mult.adder.a[14] ;
 wire \g_row[1].g_col[3].mult.adder.a[15] ;
 wire \g_row[1].g_col[3].mult.adder.a[16] ;
 wire \g_row[1].g_col[3].mult.adder.a[17] ;
 wire \g_row[1].g_col[3].mult.adder.a[18] ;
 wire \g_row[1].g_col[3].mult.adder.a[19] ;
 wire \g_row[1].g_col[3].mult.adder.a[1] ;
 wire \g_row[1].g_col[3].mult.adder.a[2] ;
 wire \g_row[1].g_col[3].mult.adder.a[3] ;
 wire \g_row[1].g_col[3].mult.adder.a[4] ;
 wire \g_row[1].g_col[3].mult.adder.a[5] ;
 wire \g_row[1].g_col[3].mult.adder.a[6] ;
 wire \g_row[1].g_col[3].mult.adder.a[7] ;
 wire \g_row[1].g_col[3].mult.adder.a[8] ;
 wire \g_row[1].g_col[3].mult.adder.a[9] ;
 wire \g_row[1].g_col[3].mult.adder.b[10] ;
 wire \g_row[1].g_col[3].mult.adder.b[11] ;
 wire \g_row[1].g_col[3].mult.adder.b[12] ;
 wire \g_row[1].g_col[3].mult.adder.b[13] ;
 wire \g_row[1].g_col[3].mult.adder.b[14] ;
 wire \g_row[1].g_col[3].mult.adder.b[15] ;
 wire \g_row[1].g_col[3].mult.adder.b[16] ;
 wire \g_row[1].g_col[3].mult.adder.b[17] ;
 wire \g_row[1].g_col[3].mult.adder.b[18] ;
 wire \g_row[1].g_col[3].mult.adder.b[19] ;
 wire \g_row[1].g_col[3].mult.adder.b[1] ;
 wire \g_row[1].g_col[3].mult.adder.b[20] ;
 wire \g_row[1].g_col[3].mult.adder.b[2] ;
 wire \g_row[1].g_col[3].mult.adder.b[3] ;
 wire \g_row[1].g_col[3].mult.adder.b[4] ;
 wire \g_row[1].g_col[3].mult.adder.b[5] ;
 wire \g_row[1].g_col[3].mult.adder.b[6] ;
 wire \g_row[1].g_col[3].mult.adder.b[7] ;
 wire \g_row[1].g_col[3].mult.adder.b[8] ;
 wire \g_row[1].g_col[3].mult.adder.b[9] ;
 wire \g_row[1].g_col[3].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[1].g_col[3].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[1].g_col[3].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[1].g_col[3].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[1].g_col[3].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[1].g_col[3].mult.sign ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[0] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[10] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[11] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[12] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[13] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[14] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[15] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[16] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[17] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[18] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[19] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[1] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[2] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[3] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[4] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[5] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[6] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[7] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[8] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t1[9] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[10] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[11] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[12] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[13] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[14] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[15] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[16] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[17] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[18] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[19] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[1] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[20] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[2] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[3] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[4] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[5] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[6] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[7] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[8] ;
 wire \g_row[1].g_col[3].mult.stage1.dadda.t2[9] ;
 wire \g_row[2].g_col[0].mult.adder.a[0] ;
 wire \g_row[2].g_col[0].mult.adder.a[10] ;
 wire \g_row[2].g_col[0].mult.adder.a[11] ;
 wire \g_row[2].g_col[0].mult.adder.a[12] ;
 wire \g_row[2].g_col[0].mult.adder.a[13] ;
 wire \g_row[2].g_col[0].mult.adder.a[14] ;
 wire \g_row[2].g_col[0].mult.adder.a[15] ;
 wire \g_row[2].g_col[0].mult.adder.a[16] ;
 wire \g_row[2].g_col[0].mult.adder.a[17] ;
 wire \g_row[2].g_col[0].mult.adder.a[18] ;
 wire \g_row[2].g_col[0].mult.adder.a[19] ;
 wire \g_row[2].g_col[0].mult.adder.a[1] ;
 wire \g_row[2].g_col[0].mult.adder.a[2] ;
 wire \g_row[2].g_col[0].mult.adder.a[3] ;
 wire \g_row[2].g_col[0].mult.adder.a[4] ;
 wire \g_row[2].g_col[0].mult.adder.a[5] ;
 wire \g_row[2].g_col[0].mult.adder.a[6] ;
 wire \g_row[2].g_col[0].mult.adder.a[7] ;
 wire \g_row[2].g_col[0].mult.adder.a[8] ;
 wire \g_row[2].g_col[0].mult.adder.a[9] ;
 wire \g_row[2].g_col[0].mult.adder.b[10] ;
 wire \g_row[2].g_col[0].mult.adder.b[11] ;
 wire \g_row[2].g_col[0].mult.adder.b[12] ;
 wire \g_row[2].g_col[0].mult.adder.b[13] ;
 wire \g_row[2].g_col[0].mult.adder.b[14] ;
 wire \g_row[2].g_col[0].mult.adder.b[15] ;
 wire \g_row[2].g_col[0].mult.adder.b[16] ;
 wire \g_row[2].g_col[0].mult.adder.b[17] ;
 wire \g_row[2].g_col[0].mult.adder.b[18] ;
 wire \g_row[2].g_col[0].mult.adder.b[19] ;
 wire \g_row[2].g_col[0].mult.adder.b[1] ;
 wire \g_row[2].g_col[0].mult.adder.b[20] ;
 wire \g_row[2].g_col[0].mult.adder.b[2] ;
 wire \g_row[2].g_col[0].mult.adder.b[3] ;
 wire \g_row[2].g_col[0].mult.adder.b[4] ;
 wire \g_row[2].g_col[0].mult.adder.b[5] ;
 wire \g_row[2].g_col[0].mult.adder.b[6] ;
 wire \g_row[2].g_col[0].mult.adder.b[7] ;
 wire \g_row[2].g_col[0].mult.adder.b[8] ;
 wire \g_row[2].g_col[0].mult.adder.b[9] ;
 wire \g_row[2].g_col[0].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[2].g_col[0].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[2].g_col[0].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[2].g_col[0].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[2].g_col[0].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[2].g_col[0].mult.sign ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[0] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[10] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[11] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[12] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[13] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[14] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[15] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[16] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[17] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[18] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[19] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[1] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[2] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[3] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[4] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[5] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[6] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[7] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[8] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t1[9] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[10] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[11] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[12] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[13] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[14] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[15] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[16] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[17] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[18] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[19] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[1] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[20] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[2] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[3] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[4] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[5] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[6] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[7] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[8] ;
 wire \g_row[2].g_col[0].mult.stage1.dadda.t2[9] ;
 wire \g_row[2].g_col[1].mult.adder.a[0] ;
 wire \g_row[2].g_col[1].mult.adder.a[10] ;
 wire \g_row[2].g_col[1].mult.adder.a[11] ;
 wire \g_row[2].g_col[1].mult.adder.a[12] ;
 wire \g_row[2].g_col[1].mult.adder.a[13] ;
 wire \g_row[2].g_col[1].mult.adder.a[14] ;
 wire \g_row[2].g_col[1].mult.adder.a[15] ;
 wire \g_row[2].g_col[1].mult.adder.a[16] ;
 wire \g_row[2].g_col[1].mult.adder.a[17] ;
 wire \g_row[2].g_col[1].mult.adder.a[18] ;
 wire \g_row[2].g_col[1].mult.adder.a[19] ;
 wire \g_row[2].g_col[1].mult.adder.a[1] ;
 wire \g_row[2].g_col[1].mult.adder.a[2] ;
 wire \g_row[2].g_col[1].mult.adder.a[3] ;
 wire \g_row[2].g_col[1].mult.adder.a[4] ;
 wire \g_row[2].g_col[1].mult.adder.a[5] ;
 wire \g_row[2].g_col[1].mult.adder.a[6] ;
 wire \g_row[2].g_col[1].mult.adder.a[7] ;
 wire \g_row[2].g_col[1].mult.adder.a[8] ;
 wire \g_row[2].g_col[1].mult.adder.a[9] ;
 wire \g_row[2].g_col[1].mult.adder.b[10] ;
 wire \g_row[2].g_col[1].mult.adder.b[11] ;
 wire \g_row[2].g_col[1].mult.adder.b[12] ;
 wire \g_row[2].g_col[1].mult.adder.b[13] ;
 wire \g_row[2].g_col[1].mult.adder.b[14] ;
 wire \g_row[2].g_col[1].mult.adder.b[15] ;
 wire \g_row[2].g_col[1].mult.adder.b[16] ;
 wire \g_row[2].g_col[1].mult.adder.b[17] ;
 wire \g_row[2].g_col[1].mult.adder.b[18] ;
 wire \g_row[2].g_col[1].mult.adder.b[19] ;
 wire \g_row[2].g_col[1].mult.adder.b[1] ;
 wire \g_row[2].g_col[1].mult.adder.b[20] ;
 wire \g_row[2].g_col[1].mult.adder.b[2] ;
 wire \g_row[2].g_col[1].mult.adder.b[3] ;
 wire \g_row[2].g_col[1].mult.adder.b[4] ;
 wire \g_row[2].g_col[1].mult.adder.b[5] ;
 wire \g_row[2].g_col[1].mult.adder.b[6] ;
 wire \g_row[2].g_col[1].mult.adder.b[7] ;
 wire \g_row[2].g_col[1].mult.adder.b[8] ;
 wire \g_row[2].g_col[1].mult.adder.b[9] ;
 wire \g_row[2].g_col[1].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[2].g_col[1].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[2].g_col[1].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[2].g_col[1].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[2].g_col[1].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[2].g_col[1].mult.sign ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[0] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[10] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[11] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[12] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[13] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[14] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[15] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[16] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[17] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[18] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[19] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[1] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[2] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[3] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[4] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[5] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[6] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[7] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[8] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t1[9] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[10] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[11] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[12] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[13] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[14] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[15] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[16] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[17] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[18] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[19] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[1] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[20] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[2] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[3] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[4] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[5] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[6] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[7] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[8] ;
 wire \g_row[2].g_col[1].mult.stage1.dadda.t2[9] ;
 wire \g_row[2].g_col[2].mult.adder.a[0] ;
 wire \g_row[2].g_col[2].mult.adder.a[10] ;
 wire \g_row[2].g_col[2].mult.adder.a[11] ;
 wire \g_row[2].g_col[2].mult.adder.a[12] ;
 wire \g_row[2].g_col[2].mult.adder.a[13] ;
 wire \g_row[2].g_col[2].mult.adder.a[14] ;
 wire \g_row[2].g_col[2].mult.adder.a[15] ;
 wire \g_row[2].g_col[2].mult.adder.a[16] ;
 wire \g_row[2].g_col[2].mult.adder.a[17] ;
 wire \g_row[2].g_col[2].mult.adder.a[18] ;
 wire \g_row[2].g_col[2].mult.adder.a[19] ;
 wire \g_row[2].g_col[2].mult.adder.a[1] ;
 wire \g_row[2].g_col[2].mult.adder.a[2] ;
 wire \g_row[2].g_col[2].mult.adder.a[3] ;
 wire \g_row[2].g_col[2].mult.adder.a[4] ;
 wire \g_row[2].g_col[2].mult.adder.a[5] ;
 wire \g_row[2].g_col[2].mult.adder.a[6] ;
 wire \g_row[2].g_col[2].mult.adder.a[7] ;
 wire \g_row[2].g_col[2].mult.adder.a[8] ;
 wire \g_row[2].g_col[2].mult.adder.a[9] ;
 wire \g_row[2].g_col[2].mult.adder.b[10] ;
 wire \g_row[2].g_col[2].mult.adder.b[11] ;
 wire \g_row[2].g_col[2].mult.adder.b[12] ;
 wire \g_row[2].g_col[2].mult.adder.b[13] ;
 wire \g_row[2].g_col[2].mult.adder.b[14] ;
 wire \g_row[2].g_col[2].mult.adder.b[15] ;
 wire \g_row[2].g_col[2].mult.adder.b[16] ;
 wire \g_row[2].g_col[2].mult.adder.b[17] ;
 wire \g_row[2].g_col[2].mult.adder.b[18] ;
 wire \g_row[2].g_col[2].mult.adder.b[19] ;
 wire \g_row[2].g_col[2].mult.adder.b[1] ;
 wire \g_row[2].g_col[2].mult.adder.b[20] ;
 wire \g_row[2].g_col[2].mult.adder.b[2] ;
 wire \g_row[2].g_col[2].mult.adder.b[3] ;
 wire \g_row[2].g_col[2].mult.adder.b[4] ;
 wire \g_row[2].g_col[2].mult.adder.b[5] ;
 wire \g_row[2].g_col[2].mult.adder.b[6] ;
 wire \g_row[2].g_col[2].mult.adder.b[7] ;
 wire \g_row[2].g_col[2].mult.adder.b[8] ;
 wire \g_row[2].g_col[2].mult.adder.b[9] ;
 wire \g_row[2].g_col[2].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[2].g_col[2].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[2].g_col[2].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[2].g_col[2].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[2].g_col[2].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[2].g_col[2].mult.sign ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[0] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[10] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[11] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[12] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[13] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[14] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[15] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[16] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[17] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[18] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[19] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[1] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[2] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[3] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[4] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[5] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[6] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[7] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[8] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t1[9] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[10] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[11] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[12] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[13] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[14] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[15] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[16] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[17] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[18] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[19] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[1] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[20] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[2] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[3] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[4] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[5] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[6] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[7] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[8] ;
 wire \g_row[2].g_col[2].mult.stage1.dadda.t2[9] ;
 wire \g_row[2].g_col[3].mult.adder.a[0] ;
 wire \g_row[2].g_col[3].mult.adder.a[10] ;
 wire \g_row[2].g_col[3].mult.adder.a[11] ;
 wire \g_row[2].g_col[3].mult.adder.a[12] ;
 wire \g_row[2].g_col[3].mult.adder.a[13] ;
 wire \g_row[2].g_col[3].mult.adder.a[14] ;
 wire \g_row[2].g_col[3].mult.adder.a[15] ;
 wire \g_row[2].g_col[3].mult.adder.a[16] ;
 wire \g_row[2].g_col[3].mult.adder.a[17] ;
 wire \g_row[2].g_col[3].mult.adder.a[18] ;
 wire \g_row[2].g_col[3].mult.adder.a[19] ;
 wire \g_row[2].g_col[3].mult.adder.a[1] ;
 wire \g_row[2].g_col[3].mult.adder.a[2] ;
 wire \g_row[2].g_col[3].mult.adder.a[3] ;
 wire \g_row[2].g_col[3].mult.adder.a[4] ;
 wire \g_row[2].g_col[3].mult.adder.a[5] ;
 wire \g_row[2].g_col[3].mult.adder.a[6] ;
 wire \g_row[2].g_col[3].mult.adder.a[7] ;
 wire \g_row[2].g_col[3].mult.adder.a[8] ;
 wire \g_row[2].g_col[3].mult.adder.a[9] ;
 wire \g_row[2].g_col[3].mult.adder.b[10] ;
 wire \g_row[2].g_col[3].mult.adder.b[11] ;
 wire \g_row[2].g_col[3].mult.adder.b[12] ;
 wire \g_row[2].g_col[3].mult.adder.b[13] ;
 wire \g_row[2].g_col[3].mult.adder.b[14] ;
 wire \g_row[2].g_col[3].mult.adder.b[15] ;
 wire \g_row[2].g_col[3].mult.adder.b[16] ;
 wire \g_row[2].g_col[3].mult.adder.b[17] ;
 wire \g_row[2].g_col[3].mult.adder.b[18] ;
 wire \g_row[2].g_col[3].mult.adder.b[19] ;
 wire \g_row[2].g_col[3].mult.adder.b[1] ;
 wire \g_row[2].g_col[3].mult.adder.b[20] ;
 wire \g_row[2].g_col[3].mult.adder.b[2] ;
 wire \g_row[2].g_col[3].mult.adder.b[3] ;
 wire \g_row[2].g_col[3].mult.adder.b[4] ;
 wire \g_row[2].g_col[3].mult.adder.b[5] ;
 wire \g_row[2].g_col[3].mult.adder.b[6] ;
 wire \g_row[2].g_col[3].mult.adder.b[7] ;
 wire \g_row[2].g_col[3].mult.adder.b[8] ;
 wire \g_row[2].g_col[3].mult.adder.b[9] ;
 wire \g_row[2].g_col[3].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[2].g_col[3].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[2].g_col[3].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[2].g_col[3].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[2].g_col[3].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[2].g_col[3].mult.sign ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[0] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[10] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[11] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[12] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[13] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[14] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[15] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[16] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[17] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[18] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[19] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[1] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[2] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[3] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[4] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[5] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[6] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[7] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[8] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t1[9] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[10] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[11] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[12] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[13] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[14] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[15] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[16] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[17] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[18] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[19] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[1] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[20] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[2] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[3] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[4] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[5] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[6] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[7] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[8] ;
 wire \g_row[2].g_col[3].mult.stage1.dadda.t2[9] ;
 wire \g_row[3].g_col[0].mult.adder.a[0] ;
 wire \g_row[3].g_col[0].mult.adder.a[10] ;
 wire \g_row[3].g_col[0].mult.adder.a[11] ;
 wire \g_row[3].g_col[0].mult.adder.a[12] ;
 wire \g_row[3].g_col[0].mult.adder.a[13] ;
 wire \g_row[3].g_col[0].mult.adder.a[14] ;
 wire \g_row[3].g_col[0].mult.adder.a[15] ;
 wire \g_row[3].g_col[0].mult.adder.a[16] ;
 wire \g_row[3].g_col[0].mult.adder.a[17] ;
 wire \g_row[3].g_col[0].mult.adder.a[18] ;
 wire \g_row[3].g_col[0].mult.adder.a[19] ;
 wire \g_row[3].g_col[0].mult.adder.a[1] ;
 wire \g_row[3].g_col[0].mult.adder.a[2] ;
 wire \g_row[3].g_col[0].mult.adder.a[3] ;
 wire \g_row[3].g_col[0].mult.adder.a[4] ;
 wire \g_row[3].g_col[0].mult.adder.a[5] ;
 wire \g_row[3].g_col[0].mult.adder.a[6] ;
 wire \g_row[3].g_col[0].mult.adder.a[7] ;
 wire \g_row[3].g_col[0].mult.adder.a[8] ;
 wire \g_row[3].g_col[0].mult.adder.a[9] ;
 wire \g_row[3].g_col[0].mult.adder.b[10] ;
 wire \g_row[3].g_col[0].mult.adder.b[11] ;
 wire \g_row[3].g_col[0].mult.adder.b[12] ;
 wire \g_row[3].g_col[0].mult.adder.b[13] ;
 wire \g_row[3].g_col[0].mult.adder.b[14] ;
 wire \g_row[3].g_col[0].mult.adder.b[15] ;
 wire \g_row[3].g_col[0].mult.adder.b[16] ;
 wire \g_row[3].g_col[0].mult.adder.b[17] ;
 wire \g_row[3].g_col[0].mult.adder.b[18] ;
 wire \g_row[3].g_col[0].mult.adder.b[19] ;
 wire \g_row[3].g_col[0].mult.adder.b[1] ;
 wire \g_row[3].g_col[0].mult.adder.b[20] ;
 wire \g_row[3].g_col[0].mult.adder.b[2] ;
 wire \g_row[3].g_col[0].mult.adder.b[3] ;
 wire \g_row[3].g_col[0].mult.adder.b[4] ;
 wire \g_row[3].g_col[0].mult.adder.b[5] ;
 wire \g_row[3].g_col[0].mult.adder.b[6] ;
 wire \g_row[3].g_col[0].mult.adder.b[7] ;
 wire \g_row[3].g_col[0].mult.adder.b[8] ;
 wire \g_row[3].g_col[0].mult.adder.b[9] ;
 wire \g_row[3].g_col[0].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[3].g_col[0].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[3].g_col[0].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[3].g_col[0].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[3].g_col[0].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[3].g_col[0].mult.sign ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[0] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[10] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[11] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[12] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[13] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[14] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[15] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[16] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[17] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[18] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[19] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[1] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[2] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[3] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[4] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[5] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[6] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[7] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[8] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t1[9] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[10] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[11] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[12] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[13] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[14] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[15] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[16] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[17] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[18] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[19] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[1] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[20] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[2] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[3] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[4] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[5] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[6] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[7] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[8] ;
 wire \g_row[3].g_col[0].mult.stage1.dadda.t2[9] ;
 wire \g_row[3].g_col[1].mult.adder.a[0] ;
 wire \g_row[3].g_col[1].mult.adder.a[10] ;
 wire \g_row[3].g_col[1].mult.adder.a[11] ;
 wire \g_row[3].g_col[1].mult.adder.a[12] ;
 wire \g_row[3].g_col[1].mult.adder.a[13] ;
 wire \g_row[3].g_col[1].mult.adder.a[14] ;
 wire \g_row[3].g_col[1].mult.adder.a[15] ;
 wire \g_row[3].g_col[1].mult.adder.a[16] ;
 wire \g_row[3].g_col[1].mult.adder.a[17] ;
 wire \g_row[3].g_col[1].mult.adder.a[18] ;
 wire \g_row[3].g_col[1].mult.adder.a[19] ;
 wire \g_row[3].g_col[1].mult.adder.a[1] ;
 wire \g_row[3].g_col[1].mult.adder.a[2] ;
 wire \g_row[3].g_col[1].mult.adder.a[3] ;
 wire \g_row[3].g_col[1].mult.adder.a[4] ;
 wire \g_row[3].g_col[1].mult.adder.a[5] ;
 wire \g_row[3].g_col[1].mult.adder.a[6] ;
 wire \g_row[3].g_col[1].mult.adder.a[7] ;
 wire \g_row[3].g_col[1].mult.adder.a[8] ;
 wire \g_row[3].g_col[1].mult.adder.a[9] ;
 wire \g_row[3].g_col[1].mult.adder.b[10] ;
 wire \g_row[3].g_col[1].mult.adder.b[11] ;
 wire \g_row[3].g_col[1].mult.adder.b[12] ;
 wire \g_row[3].g_col[1].mult.adder.b[13] ;
 wire \g_row[3].g_col[1].mult.adder.b[14] ;
 wire \g_row[3].g_col[1].mult.adder.b[15] ;
 wire \g_row[3].g_col[1].mult.adder.b[16] ;
 wire \g_row[3].g_col[1].mult.adder.b[17] ;
 wire \g_row[3].g_col[1].mult.adder.b[18] ;
 wire \g_row[3].g_col[1].mult.adder.b[19] ;
 wire \g_row[3].g_col[1].mult.adder.b[1] ;
 wire \g_row[3].g_col[1].mult.adder.b[20] ;
 wire \g_row[3].g_col[1].mult.adder.b[2] ;
 wire \g_row[3].g_col[1].mult.adder.b[3] ;
 wire \g_row[3].g_col[1].mult.adder.b[4] ;
 wire \g_row[3].g_col[1].mult.adder.b[5] ;
 wire \g_row[3].g_col[1].mult.adder.b[6] ;
 wire \g_row[3].g_col[1].mult.adder.b[7] ;
 wire \g_row[3].g_col[1].mult.adder.b[8] ;
 wire \g_row[3].g_col[1].mult.adder.b[9] ;
 wire \g_row[3].g_col[1].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[3].g_col[1].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[3].g_col[1].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[3].g_col[1].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[3].g_col[1].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[3].g_col[1].mult.sign ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[0] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[10] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[11] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[12] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[13] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[14] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[15] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[16] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[17] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[18] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[19] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[1] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[2] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[3] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[4] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[5] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[6] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[7] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[8] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t1[9] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[10] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[11] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[12] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[13] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[14] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[15] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[16] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[17] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[18] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[19] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[1] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[20] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[2] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[3] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[4] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[5] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[6] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[7] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[8] ;
 wire \g_row[3].g_col[1].mult.stage1.dadda.t2[9] ;
 wire \g_row[3].g_col[2].mult.adder.a[0] ;
 wire \g_row[3].g_col[2].mult.adder.a[10] ;
 wire \g_row[3].g_col[2].mult.adder.a[11] ;
 wire \g_row[3].g_col[2].mult.adder.a[12] ;
 wire \g_row[3].g_col[2].mult.adder.a[13] ;
 wire \g_row[3].g_col[2].mult.adder.a[14] ;
 wire \g_row[3].g_col[2].mult.adder.a[15] ;
 wire \g_row[3].g_col[2].mult.adder.a[16] ;
 wire \g_row[3].g_col[2].mult.adder.a[17] ;
 wire \g_row[3].g_col[2].mult.adder.a[18] ;
 wire \g_row[3].g_col[2].mult.adder.a[19] ;
 wire \g_row[3].g_col[2].mult.adder.a[1] ;
 wire \g_row[3].g_col[2].mult.adder.a[2] ;
 wire \g_row[3].g_col[2].mult.adder.a[3] ;
 wire \g_row[3].g_col[2].mult.adder.a[4] ;
 wire \g_row[3].g_col[2].mult.adder.a[5] ;
 wire \g_row[3].g_col[2].mult.adder.a[6] ;
 wire \g_row[3].g_col[2].mult.adder.a[7] ;
 wire \g_row[3].g_col[2].mult.adder.a[8] ;
 wire \g_row[3].g_col[2].mult.adder.a[9] ;
 wire \g_row[3].g_col[2].mult.adder.b[10] ;
 wire \g_row[3].g_col[2].mult.adder.b[11] ;
 wire \g_row[3].g_col[2].mult.adder.b[12] ;
 wire \g_row[3].g_col[2].mult.adder.b[13] ;
 wire \g_row[3].g_col[2].mult.adder.b[14] ;
 wire \g_row[3].g_col[2].mult.adder.b[15] ;
 wire \g_row[3].g_col[2].mult.adder.b[16] ;
 wire \g_row[3].g_col[2].mult.adder.b[17] ;
 wire \g_row[3].g_col[2].mult.adder.b[18] ;
 wire \g_row[3].g_col[2].mult.adder.b[19] ;
 wire \g_row[3].g_col[2].mult.adder.b[1] ;
 wire \g_row[3].g_col[2].mult.adder.b[20] ;
 wire \g_row[3].g_col[2].mult.adder.b[2] ;
 wire \g_row[3].g_col[2].mult.adder.b[3] ;
 wire \g_row[3].g_col[2].mult.adder.b[4] ;
 wire \g_row[3].g_col[2].mult.adder.b[5] ;
 wire \g_row[3].g_col[2].mult.adder.b[6] ;
 wire \g_row[3].g_col[2].mult.adder.b[7] ;
 wire \g_row[3].g_col[2].mult.adder.b[8] ;
 wire \g_row[3].g_col[2].mult.adder.b[9] ;
 wire \g_row[3].g_col[2].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[3].g_col[2].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[3].g_col[2].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[3].g_col[2].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[3].g_col[2].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[3].g_col[2].mult.sign ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[0] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[10] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[11] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[12] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[13] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[14] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[15] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[16] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[17] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[18] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[19] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[1] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[2] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[3] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[4] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[5] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[6] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[7] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[8] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t1[9] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[10] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[11] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[12] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[13] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[14] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[15] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[16] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[17] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[18] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[19] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[1] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[20] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[2] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[3] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[4] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[5] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[6] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[7] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[8] ;
 wire \g_row[3].g_col[2].mult.stage1.dadda.t2[9] ;
 wire \g_row[3].g_col[3].mult.adder.a[0] ;
 wire \g_row[3].g_col[3].mult.adder.a[10] ;
 wire \g_row[3].g_col[3].mult.adder.a[11] ;
 wire \g_row[3].g_col[3].mult.adder.a[12] ;
 wire \g_row[3].g_col[3].mult.adder.a[13] ;
 wire \g_row[3].g_col[3].mult.adder.a[14] ;
 wire \g_row[3].g_col[3].mult.adder.a[15] ;
 wire \g_row[3].g_col[3].mult.adder.a[16] ;
 wire \g_row[3].g_col[3].mult.adder.a[17] ;
 wire \g_row[3].g_col[3].mult.adder.a[18] ;
 wire \g_row[3].g_col[3].mult.adder.a[19] ;
 wire \g_row[3].g_col[3].mult.adder.a[1] ;
 wire \g_row[3].g_col[3].mult.adder.a[2] ;
 wire \g_row[3].g_col[3].mult.adder.a[3] ;
 wire \g_row[3].g_col[3].mult.adder.a[4] ;
 wire \g_row[3].g_col[3].mult.adder.a[5] ;
 wire \g_row[3].g_col[3].mult.adder.a[6] ;
 wire \g_row[3].g_col[3].mult.adder.a[7] ;
 wire \g_row[3].g_col[3].mult.adder.a[8] ;
 wire \g_row[3].g_col[3].mult.adder.a[9] ;
 wire \g_row[3].g_col[3].mult.adder.b[10] ;
 wire \g_row[3].g_col[3].mult.adder.b[11] ;
 wire \g_row[3].g_col[3].mult.adder.b[12] ;
 wire \g_row[3].g_col[3].mult.adder.b[13] ;
 wire \g_row[3].g_col[3].mult.adder.b[14] ;
 wire \g_row[3].g_col[3].mult.adder.b[15] ;
 wire \g_row[3].g_col[3].mult.adder.b[16] ;
 wire \g_row[3].g_col[3].mult.adder.b[17] ;
 wire \g_row[3].g_col[3].mult.adder.b[18] ;
 wire \g_row[3].g_col[3].mult.adder.b[19] ;
 wire \g_row[3].g_col[3].mult.adder.b[1] ;
 wire \g_row[3].g_col[3].mult.adder.b[20] ;
 wire \g_row[3].g_col[3].mult.adder.b[2] ;
 wire \g_row[3].g_col[3].mult.adder.b[3] ;
 wire \g_row[3].g_col[3].mult.adder.b[4] ;
 wire \g_row[3].g_col[3].mult.adder.b[5] ;
 wire \g_row[3].g_col[3].mult.adder.b[6] ;
 wire \g_row[3].g_col[3].mult.adder.b[7] ;
 wire \g_row[3].g_col[3].mult.adder.b[8] ;
 wire \g_row[3].g_col[3].mult.adder.b[9] ;
 wire \g_row[3].g_col[3].mult.expAdder.g_intermediate[0].fa.a ;
 wire \g_row[3].g_col[3].mult.expAdder.g_intermediate[1].fa.a ;
 wire \g_row[3].g_col[3].mult.expAdder.g_intermediate[2].fa.a ;
 wire \g_row[3].g_col[3].mult.expAdder.g_intermediate[3].fa.a ;
 wire \g_row[3].g_col[3].mult.expAdder.g_intermediate[4].fa.a ;
 wire \g_row[3].g_col[3].mult.sign ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[0] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[10] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[11] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[12] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[13] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[14] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[15] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[16] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[17] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[18] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[19] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[1] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[2] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[3] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[4] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[5] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[6] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[7] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[8] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t1[9] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[10] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[11] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[12] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[13] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[14] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[15] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[16] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[17] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[18] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[19] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[1] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[20] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[2] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[3] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[4] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[5] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[6] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[7] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[8] ;
 wire \g_row[3].g_col[3].mult.stage1.dadda.t2[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X2 _22560_ (.A(\g_reduce0[12].adder.a[12] ),
    .Z(_12154_));
 OR2_X1 _22561_ (.A1(\g_reduce0[12].adder.a[10] ),
    .A2(\g_reduce0[12].adder.a[13] ),
    .ZN(_12155_));
 OR4_X1 _22562_ (.A1(\g_reduce0[12].adder.a[11] ),
    .A2(_12154_),
    .A3(\g_reduce0[12].adder.a[14] ),
    .A4(_12155_),
    .ZN(_12156_));
 BUF_X4 _22563_ (.A(_12156_),
    .Z(_12157_));
 BUF_X2 _22564_ (.A(\g_reduce0[12].adder.b[12] ),
    .Z(_12158_));
 BUF_X2 _22565_ (.A(\g_reduce0[12].adder.b[14] ),
    .Z(_12159_));
 OR2_X1 _22566_ (.A1(\g_reduce0[12].adder.b[10] ),
    .A2(\g_reduce0[12].adder.b[13] ),
    .ZN(_12160_));
 NOR4_X4 _22567_ (.A1(\g_reduce0[12].adder.b[11] ),
    .A2(_12158_),
    .A3(_12159_),
    .A4(_12160_),
    .ZN(_12161_));
 INV_X2 _22568_ (.A(_21162_),
    .ZN(_12162_));
 CLKBUF_X3 _22569_ (.A(_21120_),
    .Z(_12163_));
 AOI21_X2 _22570_ (.A(_21119_),
    .B1(_21122_),
    .B2(_12163_),
    .ZN(_12164_));
 CLKBUF_X3 _22571_ (.A(_21123_),
    .Z(_12165_));
 NAND3_X4 _22572_ (.A1(_21162_),
    .A2(_12163_),
    .A3(_12165_),
    .ZN(_12166_));
 INV_X1 _22573_ (.A(_21128_),
    .ZN(_12167_));
 AOI21_X2 _22574_ (.A(_21125_),
    .B1(_12167_),
    .B2(_21126_),
    .ZN(_12168_));
 OAI22_X4 _22575_ (.A1(_12162_),
    .A2(_12164_),
    .B1(_12166_),
    .B2(_12168_),
    .ZN(_12169_));
 AND2_X1 _22576_ (.A1(_21132_),
    .A2(_21134_),
    .ZN(_12170_));
 BUF_X2 _22577_ (.A(_21129_),
    .Z(_12171_));
 NAND2_X1 _22578_ (.A1(_12171_),
    .A2(_21126_),
    .ZN(_12172_));
 NOR4_X1 _22579_ (.A1(_21131_),
    .A2(_12166_),
    .A3(_12170_),
    .A4(_12172_),
    .ZN(_12173_));
 AOI21_X1 _22580_ (.A(_21137_),
    .B1(_21138_),
    .B2(_21140_),
    .ZN(_12174_));
 NAND2_X1 _22581_ (.A1(_21132_),
    .A2(_21135_),
    .ZN(_12175_));
 OAI21_X2 _22582_ (.A(_12173_),
    .B1(_12174_),
    .B2(_12175_),
    .ZN(_12176_));
 AND4_X1 _22583_ (.A1(_21132_),
    .A2(_21135_),
    .A3(_21138_),
    .A4(_21141_),
    .ZN(_12177_));
 OAI22_X4 _22584_ (.A1(_21161_),
    .A2(_12169_),
    .B1(_12176_),
    .B2(_12177_),
    .ZN(_12178_));
 INV_X1 _22585_ (.A(_12178_),
    .ZN(_12179_));
 INV_X1 _22586_ (.A(_21144_),
    .ZN(_12180_));
 INV_X1 _22587_ (.A(_21146_),
    .ZN(_12181_));
 NAND2_X1 _22588_ (.A1(_21150_),
    .A2(_21153_),
    .ZN(_12182_));
 INV_X1 _22589_ (.A(\g_reduce0[12].adder.a[0] ),
    .ZN(_12183_));
 OAI21_X1 _22590_ (.A(_21156_),
    .B1(\g_reduce0[12].adder.b[0] ),
    .B2(_12183_),
    .ZN(_12184_));
 INV_X1 _22591_ (.A(_21155_),
    .ZN(_12185_));
 AOI21_X1 _22592_ (.A(_12182_),
    .B1(_12184_),
    .B2(_12185_),
    .ZN(_12186_));
 AOI21_X1 _22593_ (.A(_21149_),
    .B1(_21150_),
    .B2(_21152_),
    .ZN(_12187_));
 INV_X1 _22594_ (.A(_12187_),
    .ZN(_12188_));
 OAI21_X1 _22595_ (.A(_21147_),
    .B1(_12186_),
    .B2(_12188_),
    .ZN(_12189_));
 AOI21_X1 _22596_ (.A(_12180_),
    .B1(_12181_),
    .B2(_12189_),
    .ZN(_12190_));
 OR2_X1 _22597_ (.A1(_21143_),
    .A2(_12176_),
    .ZN(_12191_));
 OAI21_X1 _22598_ (.A(_12179_),
    .B1(_12190_),
    .B2(_12191_),
    .ZN(_12192_));
 BUF_X1 _22599_ (.A(_12192_),
    .Z(_12193_));
 OAI21_X1 _22600_ (.A(_12157_),
    .B1(_12161_),
    .B2(_12193_),
    .ZN(_12194_));
 MUX2_X2 _22601_ (.A(\g_reduce0[12].adder.a[15] ),
    .B(\g_reduce0[12].adder.b[15] ),
    .S(_12194_),
    .Z(_00038_));
 INV_X1 _22602_ (.A(_21147_),
    .ZN(_12195_));
 AND2_X1 _22603_ (.A1(_21150_),
    .A2(_21153_),
    .ZN(_12196_));
 INV_X1 _22604_ (.A(_21156_),
    .ZN(_12197_));
 INV_X1 _22605_ (.A(\g_reduce0[12].adder.b[0] ),
    .ZN(_12198_));
 AOI21_X1 _22606_ (.A(_12197_),
    .B1(_12198_),
    .B2(\g_reduce0[12].adder.a[0] ),
    .ZN(_12199_));
 OAI21_X1 _22607_ (.A(_12196_),
    .B1(_12199_),
    .B2(_21155_),
    .ZN(_12200_));
 AOI21_X1 _22608_ (.A(_12195_),
    .B1(_12200_),
    .B2(_12187_),
    .ZN(_12201_));
 OAI21_X2 _22609_ (.A(_21144_),
    .B1(_21146_),
    .B2(_12201_),
    .ZN(_12202_));
 NOR2_X1 _22610_ (.A1(_21143_),
    .A2(_12176_),
    .ZN(_12203_));
 AOI21_X4 _22611_ (.A(_12178_),
    .B1(_12202_),
    .B2(_12203_),
    .ZN(_12204_));
 CLKBUF_X3 _22612_ (.A(_12204_),
    .Z(_12205_));
 MUX2_X1 _22613_ (.A(\g_reduce0[12].adder.a[10] ),
    .B(\g_reduce0[12].adder.b[10] ),
    .S(_12205_),
    .Z(_21246_));
 INV_X1 _22614_ (.A(_12165_),
    .ZN(_12206_));
 NOR2_X1 _22615_ (.A1(\g_reduce0[12].adder.b[11] ),
    .A2(_21124_),
    .ZN(_12207_));
 INV_X1 _22616_ (.A(\g_reduce0[12].adder.b[10] ),
    .ZN(_12208_));
 OR2_X1 _22617_ (.A1(\g_reduce0[12].adder.a[10] ),
    .A2(_12208_),
    .ZN(_12209_));
 AOI21_X1 _22618_ (.A(_12207_),
    .B1(_12209_),
    .B2(_21126_),
    .ZN(_12210_));
 OAI22_X1 _22619_ (.A1(_12158_),
    .A2(_21121_),
    .B1(_12206_),
    .B2(_12210_),
    .ZN(_12211_));
 NAND2_X1 _22620_ (.A1(_12163_),
    .A2(_12211_),
    .ZN(_12212_));
 OR2_X1 _22621_ (.A1(_12163_),
    .A2(_12211_),
    .ZN(_12213_));
 AOI21_X4 _22622_ (.A(_12204_),
    .B1(_12212_),
    .B2(_12213_),
    .ZN(_12214_));
 NOR2_X1 _22623_ (.A1(\g_reduce0[12].adder.a[11] ),
    .A2(_00481_),
    .ZN(_12215_));
 NAND2_X1 _22624_ (.A1(\g_reduce0[12].adder.a[10] ),
    .A2(_12208_),
    .ZN(_12216_));
 AOI21_X1 _22625_ (.A(_12215_),
    .B1(_12216_),
    .B2(_21126_),
    .ZN(_12217_));
 OAI22_X1 _22626_ (.A1(_12154_),
    .A2(_00486_),
    .B1(_12206_),
    .B2(_12217_),
    .ZN(_12218_));
 NAND2_X1 _22627_ (.A1(_12163_),
    .A2(_12218_),
    .ZN(_12219_));
 OR2_X1 _22628_ (.A1(_12163_),
    .A2(_12218_),
    .ZN(_12220_));
 AOI21_X4 _22629_ (.A(_12192_),
    .B1(_12219_),
    .B2(_12220_),
    .ZN(_12221_));
 OR2_X2 _22630_ (.A1(_12214_),
    .A2(_12221_),
    .ZN(_12222_));
 OR2_X1 _22631_ (.A1(\g_reduce0[12].adder.b[13] ),
    .A2(_21118_),
    .ZN(_12223_));
 OAI21_X1 _22632_ (.A(_12223_),
    .B1(_21121_),
    .B2(_12158_),
    .ZN(_12224_));
 OR2_X1 _22633_ (.A1(_12165_),
    .A2(_12224_),
    .ZN(_12225_));
 OR2_X1 _22634_ (.A1(\g_reduce0[12].adder.a[13] ),
    .A2(_00489_),
    .ZN(_12226_));
 OAI21_X1 _22635_ (.A(_12226_),
    .B1(_00486_),
    .B2(_12154_),
    .ZN(_12227_));
 OR2_X1 _22636_ (.A1(_12165_),
    .A2(_12227_),
    .ZN(_12228_));
 MUX2_X2 _22637_ (.A(_12225_),
    .B(_12228_),
    .S(_12204_),
    .Z(_12229_));
 OR4_X1 _22638_ (.A1(_21158_),
    .A2(_12204_),
    .A3(_12207_),
    .A4(_12224_),
    .ZN(_12230_));
 NOR3_X1 _22639_ (.A1(_21158_),
    .A2(_12215_),
    .A3(_12227_),
    .ZN(_12231_));
 AOI21_X1 _22640_ (.A(_21162_),
    .B1(_12205_),
    .B2(_12231_),
    .ZN(_12232_));
 INV_X1 _22641_ (.A(_12163_),
    .ZN(_12233_));
 NAND2_X1 _22642_ (.A1(_12233_),
    .A2(_12223_),
    .ZN(_12234_));
 NAND2_X1 _22643_ (.A1(_12233_),
    .A2(_12226_),
    .ZN(_12235_));
 MUX2_X2 _22644_ (.A(_12234_),
    .B(_12235_),
    .S(_12204_),
    .Z(_12236_));
 NAND4_X2 _22645_ (.A1(_12229_),
    .A2(_12230_),
    .A3(_12232_),
    .A4(_12236_),
    .ZN(_12237_));
 NOR2_X1 _22646_ (.A1(_21158_),
    .A2(_12207_),
    .ZN(_12238_));
 OR2_X1 _22647_ (.A1(_12166_),
    .A2(_12238_),
    .ZN(_12239_));
 NOR2_X1 _22648_ (.A1(_21158_),
    .A2(_12215_),
    .ZN(_12240_));
 OR2_X1 _22649_ (.A1(_12166_),
    .A2(_12240_),
    .ZN(_12241_));
 MUX2_X1 _22650_ (.A(_12239_),
    .B(_12241_),
    .S(_12205_),
    .Z(_12242_));
 MUX2_X1 _22651_ (.A(_12226_),
    .B(_12223_),
    .S(_12193_),
    .Z(_12243_));
 OR3_X1 _22652_ (.A1(_12158_),
    .A2(_21121_),
    .A3(_12233_),
    .ZN(_12244_));
 OR3_X1 _22653_ (.A1(_12154_),
    .A2(_00486_),
    .A3(_12233_),
    .ZN(_12245_));
 MUX2_X1 _22654_ (.A(_12244_),
    .B(_12245_),
    .S(_12204_),
    .Z(_12246_));
 NAND4_X2 _22655_ (.A1(_21162_),
    .A2(_12242_),
    .A3(_12243_),
    .A4(_12246_),
    .ZN(_12247_));
 AND2_X2 _22656_ (.A1(_12237_),
    .A2(_12247_),
    .ZN(_12248_));
 NAND2_X2 _22657_ (.A1(_12222_),
    .A2(_12248_),
    .ZN(_12249_));
 MUX2_X1 _22658_ (.A(_00485_),
    .B(_21139_),
    .S(_12205_),
    .Z(_12250_));
 MUX2_X1 _22659_ (.A(_00484_),
    .B(_21136_),
    .S(_12205_),
    .Z(_12251_));
 INV_X2 _22660_ (.A(_12171_),
    .ZN(_12252_));
 MUX2_X1 _22661_ (.A(_12250_),
    .B(_12251_),
    .S(_12252_),
    .Z(_12253_));
 CLKBUF_X3 _22662_ (.A(_12205_),
    .Z(_12254_));
 MUX2_X1 _22663_ (.A(_00483_),
    .B(_21145_),
    .S(_12254_),
    .Z(_12255_));
 MUX2_X1 _22664_ (.A(_00482_),
    .B(_21142_),
    .S(_12254_),
    .Z(_12256_));
 MUX2_X1 _22665_ (.A(_12255_),
    .B(_12256_),
    .S(_12252_),
    .Z(_12257_));
 BUF_X2 _22666_ (.A(_21159_),
    .Z(_12258_));
 CLKBUF_X3 _22667_ (.A(_12258_),
    .Z(_12259_));
 INV_X2 _22668_ (.A(_12259_),
    .ZN(_12260_));
 MUX2_X1 _22669_ (.A(_12253_),
    .B(_12257_),
    .S(_12260_),
    .Z(_12261_));
 MUX2_X1 _22670_ (.A(_00480_),
    .B(_21151_),
    .S(_12254_),
    .Z(_12262_));
 MUX2_X1 _22671_ (.A(_00479_),
    .B(_21148_),
    .S(_12254_),
    .Z(_12263_));
 MUX2_X1 _22672_ (.A(_12262_),
    .B(_12263_),
    .S(_12252_),
    .Z(_12264_));
 MUX2_X1 _22673_ (.A(_00476_),
    .B(_21154_),
    .S(_12254_),
    .Z(_12265_));
 MUX2_X1 _22674_ (.A(_00477_),
    .B(_00478_),
    .S(_12254_),
    .Z(_12266_));
 CLKBUF_X3 _22675_ (.A(_12171_),
    .Z(_12267_));
 MUX2_X1 _22676_ (.A(_12265_),
    .B(_12266_),
    .S(_12267_),
    .Z(_12268_));
 MUX2_X1 _22677_ (.A(_12264_),
    .B(_12268_),
    .S(_12260_),
    .Z(_12269_));
 XNOR2_X2 _22678_ (.A(_12165_),
    .B(_12238_),
    .ZN(_12270_));
 INV_X1 _22679_ (.A(_12270_),
    .ZN(_12271_));
 XNOR2_X2 _22680_ (.A(_12165_),
    .B(_12240_),
    .ZN(_12272_));
 INV_X1 _22681_ (.A(_12272_),
    .ZN(_12273_));
 MUX2_X1 _22682_ (.A(_12271_),
    .B(_12273_),
    .S(_12204_),
    .Z(_12274_));
 BUF_X1 _22683_ (.A(_12274_),
    .Z(_12275_));
 MUX2_X1 _22684_ (.A(_12261_),
    .B(_12269_),
    .S(_12275_),
    .Z(_12276_));
 MUX2_X2 _22685_ (.A(_00487_),
    .B(_21130_),
    .S(_12204_),
    .Z(_12277_));
 MUX2_X1 _22686_ (.A(_00488_),
    .B(_21133_),
    .S(_12254_),
    .Z(_12278_));
 MUX2_X1 _22687_ (.A(_12277_),
    .B(_12278_),
    .S(_12267_),
    .Z(_12279_));
 MUX2_X1 _22688_ (.A(_12252_),
    .B(_12279_),
    .S(_12260_),
    .Z(_12280_));
 MUX2_X2 _22689_ (.A(_12270_),
    .B(_12272_),
    .S(_12204_),
    .Z(_12281_));
 AOI21_X4 _22690_ (.A(_12162_),
    .B1(_12229_),
    .B2(_12236_),
    .ZN(_12282_));
 AND3_X2 _22691_ (.A1(_12162_),
    .A2(_12229_),
    .A3(_12236_),
    .ZN(_12283_));
 OR4_X2 _22692_ (.A1(_12222_),
    .A2(_12281_),
    .A3(_12282_),
    .A4(_12283_),
    .ZN(_12284_));
 OAI22_X2 _22693_ (.A1(_12249_),
    .A2(_12276_),
    .B1(_12280_),
    .B2(_12284_),
    .ZN(_21223_));
 MUX2_X1 _22694_ (.A(_12262_),
    .B(_12265_),
    .S(_12267_),
    .Z(_12285_));
 NAND2_X1 _22695_ (.A1(_12260_),
    .A2(_12285_),
    .ZN(_12286_));
 MUX2_X1 _22696_ (.A(_12255_),
    .B(_12263_),
    .S(_12267_),
    .Z(_12287_));
 NAND2_X1 _22697_ (.A1(_12259_),
    .A2(_12287_),
    .ZN(_12288_));
 AND3_X1 _22698_ (.A1(_12275_),
    .A2(_12286_),
    .A3(_12288_),
    .ZN(_12289_));
 MUX2_X1 _22699_ (.A(_21133_),
    .B(_21136_),
    .S(_12171_),
    .Z(_12290_));
 OR2_X1 _22700_ (.A1(_12193_),
    .A2(_12290_),
    .ZN(_12291_));
 MUX2_X1 _22701_ (.A(_00488_),
    .B(_00484_),
    .S(_12171_),
    .Z(_12292_));
 OAI21_X1 _22702_ (.A(_12291_),
    .B1(_12292_),
    .B2(_12254_),
    .ZN(_12293_));
 NAND2_X1 _22703_ (.A1(_12259_),
    .A2(_12293_),
    .ZN(_12294_));
 MUX2_X1 _22704_ (.A(_12250_),
    .B(_12256_),
    .S(_12267_),
    .Z(_12295_));
 OAI21_X1 _22705_ (.A(_12294_),
    .B1(_12295_),
    .B2(_12259_),
    .ZN(_12296_));
 AOI21_X1 _22706_ (.A(_12289_),
    .B1(_12296_),
    .B2(_12281_),
    .ZN(_12297_));
 NOR2_X1 _22707_ (.A1(_12249_),
    .A2(_12297_),
    .ZN(_12298_));
 AOI21_X2 _22708_ (.A(_12259_),
    .B1(_12277_),
    .B2(_12267_),
    .ZN(_12299_));
 INV_X1 _22709_ (.A(_12284_),
    .ZN(_12300_));
 AOI21_X2 _22710_ (.A(_12298_),
    .B1(_12299_),
    .B2(_12300_),
    .ZN(_14064_));
 INV_X1 _22711_ (.A(_14064_),
    .ZN(_14059_));
 INV_X1 _22712_ (.A(_21223_),
    .ZN(_21226_));
 INV_X1 _22713_ (.A(_12249_),
    .ZN(_12301_));
 NAND3_X1 _22714_ (.A1(_12301_),
    .A2(_12275_),
    .A3(_12299_),
    .ZN(_21178_));
 INV_X1 _22715_ (.A(_21178_),
    .ZN(_21182_));
 OR3_X1 _22716_ (.A1(_12249_),
    .A2(_12281_),
    .A3(_12280_),
    .ZN(_21172_));
 INV_X1 _22717_ (.A(_21172_),
    .ZN(_21175_));
 NOR2_X1 _22718_ (.A1(_12252_),
    .A2(_12260_),
    .ZN(_12302_));
 MUX2_X1 _22719_ (.A(_12290_),
    .B(_12292_),
    .S(_12193_),
    .Z(_12303_));
 AOI221_X2 _22720_ (.A(_12281_),
    .B1(_12277_),
    .B2(_12302_),
    .C1(_12303_),
    .C2(_12260_),
    .ZN(_12304_));
 NAND2_X1 _22721_ (.A1(_12301_),
    .A2(_12304_),
    .ZN(_21206_));
 INV_X1 _22722_ (.A(_21206_),
    .ZN(_21210_));
 NOR2_X2 _22723_ (.A1(_12252_),
    .A2(_12259_),
    .ZN(_12305_));
 NAND2_X1 _22724_ (.A1(_12281_),
    .A2(_12305_),
    .ZN(_12306_));
 MUX2_X1 _22725_ (.A(_12253_),
    .B(_12279_),
    .S(_12259_),
    .Z(_12307_));
 OAI21_X1 _22726_ (.A(_12306_),
    .B1(_12307_),
    .B2(_12281_),
    .ZN(_12308_));
 NAND2_X1 _22727_ (.A1(_12301_),
    .A2(_12308_),
    .ZN(_21185_));
 INV_X1 _22728_ (.A(_21185_),
    .ZN(_21189_));
 MUX2_X1 _22729_ (.A(_12299_),
    .B(_12296_),
    .S(_12275_),
    .Z(_12309_));
 AND2_X1 _22730_ (.A1(_12301_),
    .A2(_12309_),
    .ZN(_21193_));
 INV_X1 _22731_ (.A(_21193_),
    .ZN(_21196_));
 MUX2_X1 _22732_ (.A(_12261_),
    .B(_12280_),
    .S(_12281_),
    .Z(_12310_));
 NOR2_X1 _22733_ (.A1(_12249_),
    .A2(_12310_),
    .ZN(_21200_));
 INV_X1 _22734_ (.A(_21200_),
    .ZN(_21203_));
 NAND2_X1 _22735_ (.A1(_12277_),
    .A2(_12302_),
    .ZN(_12311_));
 OAI21_X1 _22736_ (.A(_12311_),
    .B1(_12293_),
    .B2(_12259_),
    .ZN(_12312_));
 MUX2_X1 _22737_ (.A(_21145_),
    .B(_21139_),
    .S(_12258_),
    .Z(_12313_));
 MUX2_X1 _22738_ (.A(_21148_),
    .B(_21142_),
    .S(_12258_),
    .Z(_12314_));
 MUX2_X1 _22739_ (.A(_12313_),
    .B(_12314_),
    .S(_12267_),
    .Z(_12315_));
 MUX2_X1 _22740_ (.A(_00483_),
    .B(_00485_),
    .S(_12258_),
    .Z(_12316_));
 MUX2_X1 _22741_ (.A(_00479_),
    .B(_00482_),
    .S(_12258_),
    .Z(_12317_));
 MUX2_X1 _22742_ (.A(_12316_),
    .B(_12317_),
    .S(_12267_),
    .Z(_12318_));
 MUX2_X1 _22743_ (.A(_12315_),
    .B(_12318_),
    .S(_12193_),
    .Z(_12319_));
 MUX2_X1 _22744_ (.A(_12312_),
    .B(_12319_),
    .S(_12275_),
    .Z(_12320_));
 NOR2_X1 _22745_ (.A1(_12249_),
    .A2(_12320_),
    .ZN(_21217_));
 INV_X1 _22746_ (.A(_21217_),
    .ZN(_21220_));
 MUX2_X1 _22747_ (.A(_12257_),
    .B(_12264_),
    .S(_12260_),
    .Z(_12321_));
 MUX2_X1 _22748_ (.A(_12307_),
    .B(_12321_),
    .S(_12275_),
    .Z(_12322_));
 NOR2_X2 _22749_ (.A1(_12214_),
    .A2(_12221_),
    .ZN(_12323_));
 NAND2_X2 _22750_ (.A1(_12237_),
    .A2(_12247_),
    .ZN(_12324_));
 OAI33_X1 _22751_ (.A1(_12252_),
    .A2(_12259_),
    .A3(_12284_),
    .B1(_12322_),
    .B2(_12323_),
    .B3(_12324_),
    .ZN(_21168_));
 INV_X1 _22752_ (.A(_21168_),
    .ZN(_21213_));
 XOR2_X2 _22753_ (.A(\g_reduce0[12].adder.a[15] ),
    .B(\g_reduce0[12].adder.b[15] ),
    .Z(_12325_));
 CLKBUF_X3 _22754_ (.A(_12325_),
    .Z(_12326_));
 BUF_X2 _22755_ (.A(_21181_),
    .Z(_12327_));
 BUF_X1 _22756_ (.A(_21174_),
    .Z(_12328_));
 INV_X1 _22757_ (.A(_12328_),
    .ZN(_12329_));
 CLKBUF_X2 _22758_ (.A(_21209_),
    .Z(_12330_));
 CLKBUF_X2 _22759_ (.A(_21188_),
    .Z(_12331_));
 INV_X1 _22760_ (.A(_21194_),
    .ZN(_12332_));
 BUF_X2 _22761_ (.A(_21195_),
    .Z(_12333_));
 OAI21_X1 _22762_ (.A(_12333_),
    .B1(_21202_),
    .B2(_21201_),
    .ZN(_12334_));
 AOI21_X1 _22763_ (.A(_12331_),
    .B1(_12332_),
    .B2(_12334_),
    .ZN(_12335_));
 NOR2_X1 _22764_ (.A1(_21190_),
    .A2(_12335_),
    .ZN(_12336_));
 OR4_X1 _22765_ (.A1(_21190_),
    .A2(_21194_),
    .A3(_21201_),
    .A4(_21218_),
    .ZN(_12337_));
 INV_X1 _22766_ (.A(_21169_),
    .ZN(_12338_));
 INV_X1 _22767_ (.A(_21170_),
    .ZN(_12339_));
 AOI21_X2 _22768_ (.A(_21163_),
    .B1(_14058_),
    .B2(_21164_),
    .ZN(_12340_));
 OAI21_X4 _22769_ (.A(_12338_),
    .B1(_12339_),
    .B2(_12340_),
    .ZN(_12341_));
 BUF_X2 _22770_ (.A(_21219_),
    .Z(_12342_));
 AOI21_X2 _22771_ (.A(_12337_),
    .B1(_12341_),
    .B2(_12342_),
    .ZN(_12343_));
 NOR3_X1 _22772_ (.A1(_12330_),
    .A2(_12336_),
    .A3(_12343_),
    .ZN(_12344_));
 OAI21_X1 _22773_ (.A(_12329_),
    .B1(_12344_),
    .B2(_21211_),
    .ZN(_12345_));
 INV_X1 _22774_ (.A(_21176_),
    .ZN(_12346_));
 AOI21_X1 _22775_ (.A(_12327_),
    .B1(_12345_),
    .B2(_12346_),
    .ZN(_12347_));
 NOR2_X1 _22776_ (.A1(_21183_),
    .A2(_12347_),
    .ZN(_12348_));
 NOR2_X2 _22777_ (.A1(_12326_),
    .A2(_12348_),
    .ZN(_12349_));
 INV_X1 _22778_ (.A(_21180_),
    .ZN(_12350_));
 INV_X1 _22779_ (.A(_21208_),
    .ZN(_12351_));
 INV_X1 _22780_ (.A(_12331_),
    .ZN(_12352_));
 INV_X2 _22781_ (.A(_21197_),
    .ZN(_12353_));
 INV_X1 _22782_ (.A(_12333_),
    .ZN(_12354_));
 INV_X2 _22783_ (.A(_21202_),
    .ZN(_12355_));
 OAI21_X1 _22784_ (.A(_12354_),
    .B1(_12355_),
    .B2(_21204_),
    .ZN(_12356_));
 AOI21_X1 _22785_ (.A(_12352_),
    .B1(_12353_),
    .B2(_12356_),
    .ZN(_12357_));
 INV_X1 _22786_ (.A(_12342_),
    .ZN(_12358_));
 INV_X1 _22787_ (.A(_21214_),
    .ZN(_12359_));
 INV_X1 _22788_ (.A(_21215_),
    .ZN(_12360_));
 AOI21_X1 _22789_ (.A(_21165_),
    .B1(_14063_),
    .B2(_21166_),
    .ZN(_12361_));
 OAI21_X2 _22790_ (.A(_12359_),
    .B1(_12360_),
    .B2(_12361_),
    .ZN(_12362_));
 AND2_X1 _22791_ (.A1(_12358_),
    .A2(_12362_),
    .ZN(_12363_));
 INV_X1 _22792_ (.A(_21187_),
    .ZN(_12364_));
 INV_X1 _22793_ (.A(_21204_),
    .ZN(_12365_));
 INV_X1 _22794_ (.A(_21221_),
    .ZN(_12366_));
 NAND4_X1 _22795_ (.A1(_12353_),
    .A2(_12364_),
    .A3(_12365_),
    .A4(_12366_),
    .ZN(_12367_));
 OAI22_X1 _22796_ (.A1(_21187_),
    .A2(_12357_),
    .B1(_12363_),
    .B2(_12367_),
    .ZN(_12368_));
 INV_X1 _22797_ (.A(_12330_),
    .ZN(_12369_));
 OAI21_X1 _22798_ (.A(_12351_),
    .B1(_12368_),
    .B2(_12369_),
    .ZN(_12370_));
 AOI21_X1 _22799_ (.A(_21173_),
    .B1(_12370_),
    .B2(_12328_),
    .ZN(_12371_));
 INV_X1 _22800_ (.A(_12327_),
    .ZN(_12372_));
 OAI21_X1 _22801_ (.A(_12350_),
    .B1(_12371_),
    .B2(_12372_),
    .ZN(_12373_));
 AND2_X1 _22802_ (.A1(_12326_),
    .A2(_12373_),
    .ZN(_12374_));
 OAI211_X4 _22803_ (.A(_12275_),
    .B(_12305_),
    .C1(_12214_),
    .C2(_12221_),
    .ZN(_12375_));
 NOR4_X2 _22804_ (.A1(_12282_),
    .A2(_12283_),
    .A3(_12374_),
    .A4(_12375_),
    .ZN(_12376_));
 OR2_X2 _22805_ (.A1(_12349_),
    .A2(_12376_),
    .ZN(_12377_));
 BUF_X4 _22806_ (.A(_12377_),
    .Z(_12378_));
 XNOR2_X2 _22807_ (.A(\g_reduce0[12].adder.a[15] ),
    .B(\g_reduce0[12].adder.b[15] ),
    .ZN(_12379_));
 CLKBUF_X3 _22808_ (.A(_12379_),
    .Z(_12380_));
 NAND2_X1 _22809_ (.A1(_12329_),
    .A2(_12380_),
    .ZN(_12381_));
 OR4_X1 _22810_ (.A1(_12330_),
    .A2(_12336_),
    .A3(_12343_),
    .A4(_12381_),
    .ZN(_12382_));
 NOR3_X1 _22811_ (.A1(_21208_),
    .A2(_21173_),
    .A3(_12380_),
    .ZN(_12383_));
 NAND2_X1 _22812_ (.A1(_12353_),
    .A2(_12365_),
    .ZN(_12384_));
 AOI211_X2 _22813_ (.A(_21221_),
    .B(_12384_),
    .C1(_12362_),
    .C2(_12358_),
    .ZN(_12385_));
 AOI21_X1 _22814_ (.A(_12333_),
    .B1(_21202_),
    .B2(_12365_),
    .ZN(_12386_));
 OAI21_X1 _22815_ (.A(_12331_),
    .B1(_21197_),
    .B2(_12386_),
    .ZN(_12387_));
 OAI211_X2 _22816_ (.A(_12364_),
    .B(_12383_),
    .C1(_12385_),
    .C2(_12387_),
    .ZN(_12388_));
 NOR4_X1 _22817_ (.A1(_12330_),
    .A2(_21208_),
    .A3(_21173_),
    .A4(_12379_),
    .ZN(_12389_));
 INV_X1 _22818_ (.A(_21173_),
    .ZN(_12390_));
 MUX2_X1 _22819_ (.A(_21211_),
    .B(_12390_),
    .S(_12325_),
    .Z(_12391_));
 AOI221_X1 _22820_ (.A(_12389_),
    .B1(_12380_),
    .B2(_21176_),
    .C1(_12329_),
    .C2(_12391_),
    .ZN(_12392_));
 NAND3_X1 _22821_ (.A1(_12382_),
    .A2(_12388_),
    .A3(_12392_),
    .ZN(_12393_));
 XNOR2_X2 _22822_ (.A(_12327_),
    .B(_12393_),
    .ZN(_12394_));
 NOR2_X1 _22823_ (.A1(_12336_),
    .A2(_12343_),
    .ZN(_12395_));
 MUX2_X1 _22824_ (.A(_12395_),
    .B(_12368_),
    .S(_12325_),
    .Z(_12396_));
 XNOR2_X1 _22825_ (.A(_12330_),
    .B(_12396_),
    .ZN(_12397_));
 AOI21_X1 _22826_ (.A(_21214_),
    .B1(_14065_),
    .B2(_21215_),
    .ZN(_12398_));
 OAI21_X1 _22827_ (.A(_12366_),
    .B1(_12398_),
    .B2(_12342_),
    .ZN(_12399_));
 NOR2_X1 _22828_ (.A1(_12380_),
    .A2(_12399_),
    .ZN(_12400_));
 INV_X1 _22829_ (.A(_21218_),
    .ZN(_12401_));
 AOI21_X1 _22830_ (.A(_21169_),
    .B1(_14061_),
    .B2(_21170_),
    .ZN(_12402_));
 OAI21_X1 _22831_ (.A(_12401_),
    .B1(_12402_),
    .B2(_12358_),
    .ZN(_12403_));
 AOI21_X2 _22832_ (.A(_12400_),
    .B1(_12403_),
    .B2(_12380_),
    .ZN(_12404_));
 XNOR2_X2 _22833_ (.A(_12355_),
    .B(_12404_),
    .ZN(_12405_));
 INV_X1 _22834_ (.A(_21201_),
    .ZN(_12406_));
 AOI21_X1 _22835_ (.A(_21218_),
    .B1(_12341_),
    .B2(_12342_),
    .ZN(_12407_));
 OAI21_X1 _22836_ (.A(_12406_),
    .B1(_12407_),
    .B2(_12355_),
    .ZN(_12408_));
 OAI21_X1 _22837_ (.A(_12355_),
    .B1(_21221_),
    .B2(_12363_),
    .ZN(_12409_));
 NOR2_X1 _22838_ (.A1(_21204_),
    .A2(_12379_),
    .ZN(_12410_));
 AOI22_X2 _22839_ (.A1(_12380_),
    .A2(_12408_),
    .B1(_12409_),
    .B2(_12410_),
    .ZN(_12411_));
 XNOR2_X2 _22840_ (.A(_12333_),
    .B(_12411_),
    .ZN(_12412_));
 OR3_X1 _22841_ (.A1(_12397_),
    .A2(_12405_),
    .A3(_12412_),
    .ZN(_12413_));
 NOR2_X1 _22842_ (.A1(_12328_),
    .A2(_12380_),
    .ZN(_12414_));
 NOR2_X1 _22843_ (.A1(_12329_),
    .A2(_12380_),
    .ZN(_12415_));
 NAND3_X1 _22844_ (.A1(_12353_),
    .A2(_12364_),
    .A3(_12365_),
    .ZN(_12416_));
 AOI21_X1 _22845_ (.A(_12416_),
    .B1(_12399_),
    .B2(_12355_),
    .ZN(_12417_));
 AOI21_X1 _22846_ (.A(_12352_),
    .B1(_12353_),
    .B2(_12333_),
    .ZN(_12418_));
 OAI21_X1 _22847_ (.A(_12330_),
    .B1(_21187_),
    .B2(_12418_),
    .ZN(_12419_));
 OAI21_X1 _22848_ (.A(_12351_),
    .B1(_12417_),
    .B2(_12419_),
    .ZN(_12420_));
 MUX2_X1 _22849_ (.A(_12414_),
    .B(_12415_),
    .S(_12420_),
    .Z(_12421_));
 BUF_X4 _22850_ (.A(_12380_),
    .Z(_12422_));
 INV_X1 _22851_ (.A(_21211_),
    .ZN(_12423_));
 OAI21_X1 _22852_ (.A(_12369_),
    .B1(_21190_),
    .B2(_12352_),
    .ZN(_12424_));
 NAND2_X1 _22853_ (.A1(_12423_),
    .A2(_12424_),
    .ZN(_12425_));
 NOR3_X1 _22854_ (.A1(_21211_),
    .A2(_21190_),
    .A3(_21194_),
    .ZN(_12426_));
 AOI21_X1 _22855_ (.A(_21201_),
    .B1(_12403_),
    .B2(_21202_),
    .ZN(_12427_));
 OAI21_X2 _22856_ (.A(_12426_),
    .B1(_12427_),
    .B2(_12354_),
    .ZN(_12428_));
 AND4_X1 _22857_ (.A1(_12329_),
    .A2(_12422_),
    .A3(_12425_),
    .A4(_12428_),
    .ZN(_12429_));
 NAND2_X1 _22858_ (.A1(_12328_),
    .A2(_12380_),
    .ZN(_12430_));
 AOI21_X2 _22859_ (.A(_12430_),
    .B1(_12428_),
    .B2(_12425_),
    .ZN(_12431_));
 NOR3_X4 _22860_ (.A1(_12421_),
    .A2(_12429_),
    .A3(_12431_),
    .ZN(_12432_));
 XNOR2_X2 _22861_ (.A(_12369_),
    .B(_12396_),
    .ZN(_12433_));
 AOI21_X1 _22862_ (.A(_21204_),
    .B1(_12399_),
    .B2(_12355_),
    .ZN(_12434_));
 OAI21_X2 _22863_ (.A(_12353_),
    .B1(_12333_),
    .B2(_12434_),
    .ZN(_12435_));
 NOR2_X1 _22864_ (.A1(_21194_),
    .A2(_12325_),
    .ZN(_12436_));
 OR2_X1 _22865_ (.A1(_12354_),
    .A2(_12427_),
    .ZN(_12437_));
 AOI22_X4 _22866_ (.A1(_12326_),
    .A2(_12435_),
    .B1(_12436_),
    .B2(_12437_),
    .ZN(_12438_));
 XNOR2_X2 _22867_ (.A(_12331_),
    .B(_12438_),
    .ZN(_12439_));
 AOI21_X1 _22868_ (.A(_12432_),
    .B1(_12433_),
    .B2(_12439_),
    .ZN(_12440_));
 AOI21_X1 _22869_ (.A(_12394_),
    .B1(_12413_),
    .B2(_12440_),
    .ZN(_12441_));
 NOR2_X1 _22870_ (.A1(_21183_),
    .A2(_12326_),
    .ZN(_12442_));
 NAND3_X1 _22871_ (.A1(_12329_),
    .A2(_12425_),
    .A3(_12428_),
    .ZN(_12443_));
 AND2_X1 _22872_ (.A1(_12346_),
    .A2(_12443_),
    .ZN(_12444_));
 OAI21_X2 _22873_ (.A(_12442_),
    .B1(_12444_),
    .B2(_12327_),
    .ZN(_12445_));
 NAND2_X1 _22874_ (.A1(_12328_),
    .A2(_12420_),
    .ZN(_12446_));
 NAND3_X1 _22875_ (.A1(_12350_),
    .A2(_12390_),
    .A3(_12446_),
    .ZN(_12447_));
 AOI21_X2 _22876_ (.A(_21180_),
    .B1(_12447_),
    .B2(_12327_),
    .ZN(_12448_));
 OAI21_X4 _22877_ (.A(_12445_),
    .B1(_12448_),
    .B2(_12422_),
    .ZN(_12449_));
 NOR2_X1 _22878_ (.A1(_12441_),
    .A2(_12449_),
    .ZN(_12450_));
 INV_X1 _22879_ (.A(_12394_),
    .ZN(_12451_));
 BUF_X1 _22880_ (.A(_12397_),
    .Z(_12452_));
 NOR3_X1 _22881_ (.A1(_12452_),
    .A2(_12405_),
    .A3(_12412_),
    .ZN(_12453_));
 OR3_X1 _22882_ (.A1(_12421_),
    .A2(_12429_),
    .A3(_12431_),
    .ZN(_12454_));
 XNOR2_X2 _22883_ (.A(_12352_),
    .B(_12438_),
    .ZN(_12455_));
 OAI21_X1 _22884_ (.A(_12454_),
    .B1(_12452_),
    .B2(_12455_),
    .ZN(_12456_));
 OAI21_X1 _22885_ (.A(_12451_),
    .B1(_12453_),
    .B2(_12456_),
    .ZN(_12457_));
 AND2_X1 _22886_ (.A1(_12457_),
    .A2(_12449_),
    .ZN(_12458_));
 NOR3_X4 _22887_ (.A1(_12282_),
    .A2(_12283_),
    .A3(_12375_),
    .ZN(_12459_));
 MUX2_X1 _22888_ (.A(_12450_),
    .B(_12458_),
    .S(_12459_),
    .Z(_12460_));
 CLKBUF_X3 _22889_ (.A(_12460_),
    .Z(_12461_));
 NOR2_X1 _22890_ (.A1(_12378_),
    .A2(_12461_),
    .ZN(_12462_));
 XOR2_X1 _22891_ (.A(_14061_),
    .B(_21170_),
    .Z(_12463_));
 XOR2_X1 _22892_ (.A(_14065_),
    .B(_21215_),
    .Z(_12464_));
 MUX2_X1 _22893_ (.A(_12463_),
    .B(_12464_),
    .S(_12326_),
    .Z(_12465_));
 MUX2_X1 _22894_ (.A(_21225_),
    .B(_21227_),
    .S(_12325_),
    .Z(_12466_));
 BUF_X4 _22895_ (.A(_12466_),
    .Z(_12467_));
 NOR2_X2 _22896_ (.A1(_12465_),
    .A2(_12467_),
    .ZN(_12468_));
 NAND2_X1 _22897_ (.A1(_12422_),
    .A2(_12468_),
    .ZN(_12469_));
 NOR3_X1 _22898_ (.A1(_12214_),
    .A2(_12221_),
    .A3(_12469_),
    .ZN(_12470_));
 NAND4_X2 _22899_ (.A1(_12237_),
    .A2(_12247_),
    .A3(_12304_),
    .A4(_12470_),
    .ZN(_12471_));
 NAND2_X1 _22900_ (.A1(_12326_),
    .A2(_12468_),
    .ZN(_12472_));
 OAI21_X4 _22901_ (.A(_12471_),
    .B1(_12472_),
    .B2(_12248_),
    .ZN(_12473_));
 NAND2_X1 _22902_ (.A1(_12171_),
    .A2(_12259_),
    .ZN(_12474_));
 MUX2_X1 _22903_ (.A(_00478_),
    .B(_21151_),
    .S(_12258_),
    .Z(_12475_));
 OAI22_X1 _22904_ (.A1(_21154_),
    .A2(_12474_),
    .B1(_12475_),
    .B2(_12267_),
    .ZN(_12476_));
 OR3_X1 _22905_ (.A1(_12193_),
    .A2(_12272_),
    .A3(_12476_),
    .ZN(_12477_));
 NAND3_X1 _22906_ (.A1(_12205_),
    .A2(_12272_),
    .A3(_12315_),
    .ZN(_12478_));
 NAND3_X1 _22907_ (.A1(_12193_),
    .A2(_12270_),
    .A3(_12318_),
    .ZN(_12479_));
 MUX2_X1 _22908_ (.A(_00477_),
    .B(_00480_),
    .S(_12258_),
    .Z(_12480_));
 OAI22_X1 _22909_ (.A1(_00476_),
    .A2(_12474_),
    .B1(_12480_),
    .B2(_12267_),
    .ZN(_12481_));
 OR3_X1 _22910_ (.A1(_12204_),
    .A2(_12270_),
    .A3(_12481_),
    .ZN(_12482_));
 NAND4_X4 _22911_ (.A1(_12477_),
    .A2(_12478_),
    .A3(_12479_),
    .A4(_12482_),
    .ZN(_12483_));
 NAND4_X2 _22912_ (.A1(_12222_),
    .A2(_12326_),
    .A3(_12468_),
    .A4(_12483_),
    .ZN(_12484_));
 OR3_X1 _22913_ (.A1(_12222_),
    .A2(_12304_),
    .A3(_12472_),
    .ZN(_12485_));
 OR3_X1 _22914_ (.A1(_12323_),
    .A2(_12483_),
    .A3(_12469_),
    .ZN(_12486_));
 OAI211_X4 _22915_ (.A(_12484_),
    .B(_12485_),
    .C1(_12324_),
    .C2(_12486_),
    .ZN(_12487_));
 BUF_X2 _22916_ (.A(_12394_),
    .Z(_12488_));
 NOR2_X1 _22917_ (.A1(_12422_),
    .A2(_12362_),
    .ZN(_12489_));
 AOI21_X4 _22918_ (.A(_12489_),
    .B1(_12341_),
    .B2(_12422_),
    .ZN(_12490_));
 XNOR2_X2 _22919_ (.A(_12358_),
    .B(_12490_),
    .ZN(_12491_));
 AND2_X1 _22920_ (.A1(_14062_),
    .A2(_12422_),
    .ZN(_12492_));
 AND2_X1 _22921_ (.A1(_14066_),
    .A2(_12326_),
    .ZN(_12493_));
 OR2_X2 _22922_ (.A1(_12492_),
    .A2(_12493_),
    .ZN(_12494_));
 OAI21_X1 _22923_ (.A(_12491_),
    .B1(_12494_),
    .B2(_12465_),
    .ZN(_12495_));
 NOR2_X1 _22924_ (.A1(_12488_),
    .A2(_12495_),
    .ZN(_12496_));
 AOI21_X2 _22925_ (.A(_12452_),
    .B1(_12455_),
    .B2(_12412_),
    .ZN(_12497_));
 OAI21_X2 _22926_ (.A(_12496_),
    .B1(_12497_),
    .B2(_12432_),
    .ZN(_12498_));
 NOR4_X4 _22927_ (.A1(_12377_),
    .A2(_12473_),
    .A3(_12487_),
    .A4(_12498_),
    .ZN(_12499_));
 NOR2_X4 _22928_ (.A1(_12462_),
    .A2(_12499_),
    .ZN(_21229_));
 INV_X1 _22929_ (.A(_21229_),
    .ZN(_21231_));
 INV_X1 _22930_ (.A(_21234_),
    .ZN(_12500_));
 OR2_X1 _22931_ (.A1(_12394_),
    .A2(_12432_),
    .ZN(_12501_));
 NOR3_X2 _22932_ (.A1(_12452_),
    .A2(_12439_),
    .A3(_12501_),
    .ZN(_12502_));
 CLKBUF_X3 _22933_ (.A(_12465_),
    .Z(_12503_));
 XNOR2_X2 _22934_ (.A(_12342_),
    .B(_12490_),
    .ZN(_12504_));
 OR2_X2 _22935_ (.A1(_12503_),
    .A2(_12504_),
    .ZN(_12505_));
 INV_X1 _22936_ (.A(_12412_),
    .ZN(_12506_));
 NAND2_X1 _22937_ (.A1(_12405_),
    .A2(_12506_),
    .ZN(_12507_));
 OAI21_X2 _22938_ (.A(_12502_),
    .B1(_12505_),
    .B2(_12507_),
    .ZN(_12508_));
 AND3_X1 _22939_ (.A1(_12326_),
    .A2(_12373_),
    .A3(_12447_),
    .ZN(_12509_));
 NAND4_X1 _22940_ (.A1(_12222_),
    .A2(_12275_),
    .A3(_12305_),
    .A4(_12509_),
    .ZN(_12510_));
 OAI33_X1 _22941_ (.A1(_12349_),
    .A2(_12459_),
    .A3(_12449_),
    .B1(_12510_),
    .B2(_12282_),
    .B3(_12283_),
    .ZN(_12511_));
 BUF_X4 _22942_ (.A(_12511_),
    .Z(_12512_));
 AOI21_X4 _22943_ (.A(_12500_),
    .B1(_12508_),
    .B2(_12512_),
    .ZN(_12513_));
 AND3_X2 _22944_ (.A1(_12500_),
    .A2(_12508_),
    .A3(_12512_),
    .ZN(_12514_));
 NOR2_X4 _22945_ (.A1(_12513_),
    .A2(_12514_),
    .ZN(_12515_));
 INV_X1 _22946_ (.A(_12515_),
    .ZN(_21255_));
 NAND3_X1 _22947_ (.A1(_12323_),
    .A2(_12304_),
    .A3(_12422_),
    .ZN(_12516_));
 MUX2_X2 _22948_ (.A(_12422_),
    .B(_12516_),
    .S(_12248_),
    .Z(_12517_));
 NOR3_X1 _22949_ (.A1(_12222_),
    .A2(_12304_),
    .A3(_12422_),
    .ZN(_12518_));
 NOR2_X1 _22950_ (.A1(_12323_),
    .A2(_12422_),
    .ZN(_12519_));
 NOR3_X1 _22951_ (.A1(_12323_),
    .A2(_12326_),
    .A3(_12483_),
    .ZN(_12520_));
 AOI221_X2 _22952_ (.A(_12518_),
    .B1(_12519_),
    .B2(_12483_),
    .C1(_12520_),
    .C2(_12248_),
    .ZN(_12521_));
 NAND2_X2 _22953_ (.A1(_12517_),
    .A2(_12521_),
    .ZN(_12522_));
 NOR3_X1 _22954_ (.A1(_12349_),
    .A2(_12459_),
    .A3(_12449_),
    .ZN(_12523_));
 AOI21_X2 _22955_ (.A(_12523_),
    .B1(_12509_),
    .B2(_12459_),
    .ZN(_12524_));
 NAND2_X1 _22956_ (.A1(_12522_),
    .A2(_12524_),
    .ZN(_12525_));
 BUF_X4 _22957_ (.A(_12498_),
    .Z(_12526_));
 INV_X1 _22958_ (.A(_12526_),
    .ZN(_12527_));
 OR2_X1 _22959_ (.A1(_12441_),
    .A2(_12449_),
    .ZN(_12528_));
 NAND2_X1 _22960_ (.A1(_12457_),
    .A2(_12449_),
    .ZN(_12529_));
 MUX2_X1 _22961_ (.A(_12528_),
    .B(_12529_),
    .S(_12459_),
    .Z(_12530_));
 BUF_X4 _22962_ (.A(_12530_),
    .Z(_12531_));
 OAI211_X4 _22963_ (.A(_12517_),
    .B(_12521_),
    .C1(_12527_),
    .C2(_12531_),
    .ZN(_12532_));
 BUF_X2 _22964_ (.A(_14068_),
    .Z(_12533_));
 INV_X1 _22965_ (.A(_12533_),
    .ZN(_12534_));
 NOR2_X1 _22966_ (.A1(_12534_),
    .A2(_12378_),
    .ZN(_12535_));
 OAI211_X2 _22967_ (.A(_12532_),
    .B(_12535_),
    .C1(_12513_),
    .C2(_12514_),
    .ZN(_12536_));
 NOR2_X2 _22968_ (.A1(_12349_),
    .A2(_12376_),
    .ZN(_12537_));
 INV_X1 _22969_ (.A(_12405_),
    .ZN(_12538_));
 NOR2_X1 _22970_ (.A1(_12538_),
    .A2(_12412_),
    .ZN(_12539_));
 NOR2_X2 _22971_ (.A1(_12492_),
    .A2(_12493_),
    .ZN(_12540_));
 NOR2_X1 _22972_ (.A1(_12467_),
    .A2(_12540_),
    .ZN(_12541_));
 OAI21_X1 _22973_ (.A(_12539_),
    .B1(_12541_),
    .B2(_12505_),
    .ZN(_12542_));
 NAND2_X1 _22974_ (.A1(_12455_),
    .A2(_12495_),
    .ZN(_12543_));
 AOI21_X1 _22975_ (.A(_12432_),
    .B1(_12497_),
    .B2(_12543_),
    .ZN(_12544_));
 OAI33_X1 _22976_ (.A1(_12538_),
    .A2(_12412_),
    .A3(_12505_),
    .B1(_12542_),
    .B2(_12544_),
    .B3(_12488_),
    .ZN(_12545_));
 NAND2_X1 _22977_ (.A1(_12502_),
    .A2(_12545_),
    .ZN(_12546_));
 NAND3_X4 _22978_ (.A1(_12537_),
    .A2(_12512_),
    .A3(_12546_),
    .ZN(_12547_));
 OAI21_X1 _22979_ (.A(_12525_),
    .B1(_12536_),
    .B2(_12547_),
    .ZN(_12548_));
 CLKBUF_X3 _22980_ (.A(_21230_),
    .Z(_12549_));
 CLKBUF_X3 _22981_ (.A(_12524_),
    .Z(_12550_));
 NAND2_X1 _22982_ (.A1(_12549_),
    .A2(_12550_),
    .ZN(_12551_));
 MUX2_X1 _22983_ (.A(_12467_),
    .B(_12548_),
    .S(_12551_),
    .Z(_12552_));
 INV_X1 _22984_ (.A(_12467_),
    .ZN(_12553_));
 INV_X1 _22985_ (.A(_21230_),
    .ZN(_12554_));
 CLKBUF_X3 _22986_ (.A(_12554_),
    .Z(_12555_));
 AOI21_X1 _22987_ (.A(_12512_),
    .B1(_12553_),
    .B2(_12555_),
    .ZN(_12556_));
 NOR2_X4 _22988_ (.A1(_12515_),
    .A2(_12547_),
    .ZN(_12557_));
 BUF_X4 _22989_ (.A(_12534_),
    .Z(_12558_));
 NOR3_X2 _22990_ (.A1(_12473_),
    .A2(_12487_),
    .A3(_12526_),
    .ZN(_12559_));
 OAI22_X4 _22991_ (.A1(_12558_),
    .A2(_12467_),
    .B1(_12559_),
    .B2(_12531_),
    .ZN(_12560_));
 BUF_X4 _22992_ (.A(_12533_),
    .Z(_12561_));
 NOR2_X1 _22993_ (.A1(_12468_),
    .A2(_12526_),
    .ZN(_12562_));
 NOR2_X1 _22994_ (.A1(_12531_),
    .A2(_12562_),
    .ZN(_12563_));
 NAND3_X2 _22995_ (.A1(_12561_),
    .A2(_12522_),
    .A3(_12563_),
    .ZN(_12564_));
 AOI21_X4 _22996_ (.A(_12378_),
    .B1(_12560_),
    .B2(_12564_),
    .ZN(_12565_));
 AOI21_X2 _22997_ (.A(_12556_),
    .B1(_12557_),
    .B2(_12565_),
    .ZN(_12566_));
 NOR2_X1 _22998_ (.A1(_12555_),
    .A2(_12512_),
    .ZN(_12567_));
 AOI21_X1 _22999_ (.A(_12566_),
    .B1(_12567_),
    .B2(_12494_),
    .ZN(_12568_));
 AND2_X1 _23000_ (.A1(_12552_),
    .A2(_12568_),
    .ZN(_21236_));
 NOR4_X4 _23001_ (.A1(\g_reduce0[12].adder.a[11] ),
    .A2(_12154_),
    .A3(\g_reduce0[12].adder.a[14] ),
    .A4(_12155_),
    .ZN(_12569_));
 CLKBUF_X3 _23002_ (.A(_12537_),
    .Z(_12570_));
 NOR2_X1 _23003_ (.A1(_12549_),
    .A2(_12570_),
    .ZN(_12571_));
 BUF_X4 _23004_ (.A(_12515_),
    .Z(_12572_));
 XNOR2_X2 _23005_ (.A(_12459_),
    .B(_12449_),
    .ZN(_12573_));
 AOI21_X1 _23006_ (.A(_12452_),
    .B1(_12573_),
    .B2(_12488_),
    .ZN(_12574_));
 XOR2_X2 _23007_ (.A(_12459_),
    .B(_12449_),
    .Z(_12575_));
 AOI21_X1 _23008_ (.A(_12439_),
    .B1(_12432_),
    .B2(_12451_),
    .ZN(_12576_));
 INV_X1 _23009_ (.A(_12576_),
    .ZN(_12577_));
 OAI221_X2 _23010_ (.A(_12570_),
    .B1(_12452_),
    .B2(_12439_),
    .C1(_12575_),
    .C2(_12577_),
    .ZN(_12578_));
 NOR3_X1 _23011_ (.A1(_12558_),
    .A2(_12574_),
    .A3(_12578_),
    .ZN(_12579_));
 NAND2_X1 _23012_ (.A1(_12558_),
    .A2(_12570_),
    .ZN(_12580_));
 NAND2_X1 _23013_ (.A1(_12538_),
    .A2(_12461_),
    .ZN(_12581_));
 NAND2_X1 _23014_ (.A1(_12412_),
    .A2(_12531_),
    .ZN(_12582_));
 AOI21_X1 _23015_ (.A(_12580_),
    .B1(_12581_),
    .B2(_12582_),
    .ZN(_12583_));
 OR2_X1 _23016_ (.A1(_12579_),
    .A2(_12583_),
    .ZN(_12584_));
 NAND2_X1 _23017_ (.A1(_12572_),
    .A2(_12584_),
    .ZN(_12585_));
 OAI21_X1 _23018_ (.A(_12488_),
    .B1(_12432_),
    .B2(_12575_),
    .ZN(_12586_));
 NOR2_X1 _23019_ (.A1(_12378_),
    .A2(_12586_),
    .ZN(_12587_));
 NAND3_X1 _23020_ (.A1(_12558_),
    .A2(_21255_),
    .A3(_12587_),
    .ZN(_12588_));
 AOI21_X1 _23021_ (.A(_12547_),
    .B1(_12585_),
    .B2(_12588_),
    .ZN(_12589_));
 NAND2_X1 _23022_ (.A1(_12502_),
    .A2(_12539_),
    .ZN(_12590_));
 INV_X1 _23023_ (.A(_12590_),
    .ZN(_12591_));
 OAI21_X1 _23024_ (.A(_12505_),
    .B1(_12544_),
    .B2(_12488_),
    .ZN(_12592_));
 NAND3_X2 _23025_ (.A1(_12512_),
    .A2(_12591_),
    .A3(_12592_),
    .ZN(_12593_));
 OAI21_X1 _23026_ (.A(_12540_),
    .B1(_12559_),
    .B2(_12531_),
    .ZN(_12594_));
 NAND2_X2 _23027_ (.A1(_12467_),
    .A2(_12526_),
    .ZN(_12595_));
 OAI21_X2 _23028_ (.A(_12594_),
    .B1(_12595_),
    .B2(_12531_),
    .ZN(_12596_));
 NOR2_X2 _23029_ (.A1(_12561_),
    .A2(_12572_),
    .ZN(_12597_));
 AND2_X1 _23030_ (.A1(_12503_),
    .A2(_12526_),
    .ZN(_12598_));
 MUX2_X1 _23031_ (.A(_12504_),
    .B(_12598_),
    .S(_12461_),
    .Z(_12599_));
 MUX2_X1 _23032_ (.A(_12532_),
    .B(_12599_),
    .S(_21255_),
    .Z(_12600_));
 AOI22_X4 _23033_ (.A1(_12596_),
    .A2(_12597_),
    .B1(_12600_),
    .B2(_12561_),
    .ZN(_12601_));
 NOR2_X1 _23034_ (.A1(_12593_),
    .A2(_12601_),
    .ZN(_12602_));
 OR3_X2 _23035_ (.A1(_12571_),
    .A2(_12589_),
    .A3(_12602_),
    .ZN(_12603_));
 INV_X1 _23036_ (.A(_21232_),
    .ZN(_12604_));
 NAND2_X2 _23037_ (.A1(_12570_),
    .A2(_12593_),
    .ZN(_12605_));
 NOR3_X1 _23038_ (.A1(_12604_),
    .A2(_12572_),
    .A3(_12605_),
    .ZN(_12606_));
 OAI21_X1 _23039_ (.A(_12552_),
    .B1(_12606_),
    .B2(_12550_),
    .ZN(_12607_));
 MUX2_X1 _23040_ (.A(_12607_),
    .B(_12552_),
    .S(_12568_),
    .Z(_12608_));
 OR3_X1 _23041_ (.A1(_12161_),
    .A2(_12603_),
    .A3(_12608_),
    .ZN(_12609_));
 OR4_X1 _23042_ (.A1(\g_reduce0[12].adder.b[11] ),
    .A2(_12158_),
    .A3(_12159_),
    .A4(_12160_),
    .ZN(_12610_));
 CLKBUF_X3 _23043_ (.A(_12610_),
    .Z(_12611_));
 NAND3_X1 _23044_ (.A1(_21239_),
    .A2(_12611_),
    .A3(_12603_),
    .ZN(_12612_));
 NAND2_X1 _23045_ (.A1(_12503_),
    .A2(_12550_),
    .ZN(_12613_));
 OAI22_X4 _23046_ (.A1(_12494_),
    .A2(_12526_),
    .B1(_12595_),
    .B2(_12531_),
    .ZN(_12614_));
 OAI21_X1 _23047_ (.A(_12533_),
    .B1(_12461_),
    .B2(_12494_),
    .ZN(_12615_));
 OAI221_X2 _23048_ (.A(_12570_),
    .B1(_12614_),
    .B2(_12615_),
    .C1(_12532_),
    .C2(_12533_),
    .ZN(_12616_));
 INV_X1 _23049_ (.A(_12616_),
    .ZN(_12617_));
 AOI22_X2 _23050_ (.A1(_12540_),
    .A2(_12550_),
    .B1(_12557_),
    .B2(_12617_),
    .ZN(_12618_));
 OR3_X2 _23051_ (.A1(_12513_),
    .A2(_12514_),
    .A3(_12547_),
    .ZN(_12619_));
 OAI22_X1 _23052_ (.A1(_12491_),
    .A2(_12551_),
    .B1(_12619_),
    .B2(_12604_),
    .ZN(_12620_));
 OAI211_X2 _23053_ (.A(_12461_),
    .B(_12522_),
    .C1(_12526_),
    .C2(_12468_),
    .ZN(_12621_));
 NAND4_X1 _23054_ (.A1(_12461_),
    .A2(_12517_),
    .A3(_12521_),
    .A4(_12526_),
    .ZN(_12622_));
 AOI21_X2 _23055_ (.A(_12561_),
    .B1(_12467_),
    .B2(_12622_),
    .ZN(_12623_));
 NAND2_X1 _23056_ (.A1(_12570_),
    .A2(_12531_),
    .ZN(_12624_));
 OR4_X2 _23057_ (.A1(_12378_),
    .A2(_12473_),
    .A3(_12487_),
    .A4(_12526_),
    .ZN(_12625_));
 NAND3_X2 _23058_ (.A1(_12540_),
    .A2(_12624_),
    .A3(_12625_),
    .ZN(_12626_));
 AOI21_X2 _23059_ (.A(_12378_),
    .B1(_12461_),
    .B2(_12526_),
    .ZN(_12627_));
 AOI21_X2 _23060_ (.A(_12558_),
    .B1(_12503_),
    .B2(_12627_),
    .ZN(_12628_));
 AOI22_X4 _23061_ (.A1(_12621_),
    .A2(_12623_),
    .B1(_12626_),
    .B2(_12628_),
    .ZN(_12629_));
 AOI21_X1 _23062_ (.A(_12620_),
    .B1(_12629_),
    .B2(_12557_),
    .ZN(_12630_));
 NOR2_X1 _23063_ (.A1(_12575_),
    .A2(_12605_),
    .ZN(_12631_));
 NAND2_X1 _23064_ (.A1(_12503_),
    .A2(_12631_),
    .ZN(_12632_));
 NOR2_X2 _23065_ (.A1(_12378_),
    .A2(_12572_),
    .ZN(_12633_));
 AOI22_X4 _23066_ (.A1(_21232_),
    .A2(_12572_),
    .B1(_12633_),
    .B2(_12629_),
    .ZN(_12634_));
 OAI221_X2 _23067_ (.A(_12613_),
    .B1(_12618_),
    .B2(_12630_),
    .C1(_12632_),
    .C2(_12634_),
    .ZN(_12635_));
 NAND2_X1 _23068_ (.A1(_12533_),
    .A2(_12405_),
    .ZN(_12636_));
 AOI21_X1 _23069_ (.A(_12636_),
    .B1(_12625_),
    .B2(_12624_),
    .ZN(_12637_));
 NOR2_X1 _23070_ (.A1(_12534_),
    .A2(_12504_),
    .ZN(_12638_));
 AOI21_X1 _23071_ (.A(_12533_),
    .B1(_12503_),
    .B2(_12627_),
    .ZN(_12639_));
 AOI221_X2 _23072_ (.A(_12637_),
    .B1(_12638_),
    .B2(_21229_),
    .C1(_12639_),
    .C2(_12626_),
    .ZN(_12640_));
 AOI22_X4 _23073_ (.A1(_12572_),
    .A2(_12565_),
    .B1(_12640_),
    .B2(_12633_),
    .ZN(_12641_));
 NOR2_X1 _23074_ (.A1(_12549_),
    .A2(_12405_),
    .ZN(_12642_));
 AOI21_X2 _23075_ (.A(_12642_),
    .B1(_12412_),
    .B2(_12549_),
    .ZN(_12643_));
 BUF_X4 _23076_ (.A(_12512_),
    .Z(_12644_));
 OAI22_X4 _23077_ (.A1(_12547_),
    .A2(_12641_),
    .B1(_12643_),
    .B2(_12644_),
    .ZN(_12645_));
 MUX2_X1 _23078_ (.A(_12405_),
    .B(_12491_),
    .S(_12555_),
    .Z(_12646_));
 OAI22_X4 _23079_ (.A1(_12547_),
    .A2(_12601_),
    .B1(_12646_),
    .B2(_12644_),
    .ZN(_12647_));
 OAI33_X1 _23080_ (.A1(_12492_),
    .A2(_12493_),
    .A3(_12512_),
    .B1(_12515_),
    .B2(_12547_),
    .B3(_12616_),
    .ZN(_12648_));
 NAND3_X1 _23081_ (.A1(_12551_),
    .A2(_12548_),
    .A3(_12648_),
    .ZN(_12649_));
 NAND4_X1 _23082_ (.A1(_12503_),
    .A2(_12467_),
    .A3(_12504_),
    .A4(_12567_),
    .ZN(_12650_));
 AOI221_X1 _23083_ (.A(_12566_),
    .B1(_12649_),
    .B2(_12650_),
    .C1(_12567_),
    .C2(_12494_),
    .ZN(_12651_));
 NAND4_X4 _23084_ (.A1(_12635_),
    .A2(_12645_),
    .A3(_12647_),
    .A4(_12651_),
    .ZN(_12652_));
 NOR2_X1 _23085_ (.A1(_12561_),
    .A2(_12405_),
    .ZN(_12653_));
 NOR2_X1 _23086_ (.A1(_12558_),
    .A2(_12455_),
    .ZN(_12654_));
 OAI22_X2 _23087_ (.A1(_12462_),
    .A2(_12499_),
    .B1(_12653_),
    .B2(_12654_),
    .ZN(_12655_));
 NOR2_X1 _23088_ (.A1(_12561_),
    .A2(_12491_),
    .ZN(_12656_));
 NOR2_X1 _23089_ (.A1(_12534_),
    .A2(_12506_),
    .ZN(_12657_));
 OAI221_X2 _23090_ (.A(_12625_),
    .B1(_12656_),
    .B2(_12657_),
    .C1(_12461_),
    .C2(_12378_),
    .ZN(_12658_));
 AOI21_X1 _23091_ (.A(_12619_),
    .B1(_12655_),
    .B2(_12658_),
    .ZN(_12659_));
 OAI21_X1 _23092_ (.A(_12561_),
    .B1(_12488_),
    .B2(_12575_),
    .ZN(_12660_));
 AOI21_X1 _23093_ (.A(_12433_),
    .B1(_12575_),
    .B2(_12570_),
    .ZN(_12661_));
 AOI21_X1 _23094_ (.A(_12378_),
    .B1(_12488_),
    .B2(_12573_),
    .ZN(_12662_));
 OAI22_X1 _23095_ (.A1(_12432_),
    .A2(_12661_),
    .B1(_12662_),
    .B2(_12452_),
    .ZN(_12663_));
 OAI21_X1 _23096_ (.A(_12660_),
    .B1(_12663_),
    .B2(_12561_),
    .ZN(_12664_));
 AOI21_X1 _23097_ (.A(_12659_),
    .B1(_12664_),
    .B2(_12557_),
    .ZN(_12665_));
 MUX2_X1 _23098_ (.A(_12570_),
    .B(_12573_),
    .S(_12555_),
    .Z(_12666_));
 INV_X1 _23099_ (.A(_12605_),
    .ZN(_21258_));
 OAI211_X2 _23100_ (.A(_12665_),
    .B(_12666_),
    .C1(_21258_),
    .C2(_12634_),
    .ZN(_12667_));
 NAND3_X1 _23101_ (.A1(_12549_),
    .A2(_12570_),
    .A3(_12575_),
    .ZN(_12668_));
 NAND3_X1 _23102_ (.A1(_12555_),
    .A2(_12378_),
    .A3(_12573_),
    .ZN(_12669_));
 NAND3_X2 _23103_ (.A1(_12667_),
    .A2(_12668_),
    .A3(_12669_),
    .ZN(_12670_));
 OAI22_X1 _23104_ (.A1(_12549_),
    .A2(_12488_),
    .B1(_12575_),
    .B2(_12571_),
    .ZN(_12671_));
 NOR2_X1 _23105_ (.A1(_12593_),
    .A2(_12616_),
    .ZN(_12672_));
 NOR2_X1 _23106_ (.A1(_12574_),
    .A2(_12578_),
    .ZN(_12673_));
 MUX2_X1 _23107_ (.A(_12587_),
    .B(_12673_),
    .S(_12558_),
    .Z(_12674_));
 NOR3_X1 _23108_ (.A1(_12572_),
    .A2(_12672_),
    .A3(_12674_),
    .ZN(_12675_));
 NAND2_X1 _23109_ (.A1(_12582_),
    .A2(_12581_),
    .ZN(_12676_));
 MUX2_X1 _23110_ (.A(_12599_),
    .B(_12676_),
    .S(_12561_),
    .Z(_12677_));
 NOR2_X1 _23111_ (.A1(_21255_),
    .A2(_12677_),
    .ZN(_12678_));
 OR3_X1 _23112_ (.A1(_12550_),
    .A2(_12675_),
    .A3(_12678_),
    .ZN(_12679_));
 AND2_X2 _23113_ (.A1(_12671_),
    .A2(_12679_),
    .ZN(_12680_));
 MUX2_X1 _23114_ (.A(_12452_),
    .B(_12439_),
    .S(_12554_),
    .Z(_12681_));
 NAND2_X1 _23115_ (.A1(_12524_),
    .A2(_12681_),
    .ZN(_12682_));
 OAI211_X2 _23116_ (.A(_21232_),
    .B(_12512_),
    .C1(_12513_),
    .C2(_12514_),
    .ZN(_12683_));
 OAI21_X1 _23117_ (.A(_12682_),
    .B1(_12683_),
    .B2(_21258_),
    .ZN(_12684_));
 OR3_X1 _23118_ (.A1(_12524_),
    .A2(_12513_),
    .A3(_12514_),
    .ZN(_12685_));
 NAND3_X1 _23119_ (.A1(_12500_),
    .A2(_12524_),
    .A3(_12681_),
    .ZN(_12686_));
 OAI21_X1 _23120_ (.A(_12467_),
    .B1(_12462_),
    .B2(_12499_),
    .ZN(_12687_));
 OAI21_X1 _23121_ (.A(_12570_),
    .B1(_12531_),
    .B2(_12562_),
    .ZN(_12688_));
 AOI21_X1 _23122_ (.A(_12533_),
    .B1(_12522_),
    .B2(_12688_),
    .ZN(_12689_));
 AOI221_X2 _23123_ (.A(_12605_),
    .B1(_12685_),
    .B2(_12686_),
    .C1(_12687_),
    .C2(_12689_),
    .ZN(_12690_));
 NAND2_X1 _23124_ (.A1(_12626_),
    .A2(_12628_),
    .ZN(_12691_));
 NAND2_X1 _23125_ (.A1(_12655_),
    .A2(_12658_),
    .ZN(_12692_));
 NOR2_X1 _23126_ (.A1(_12550_),
    .A2(_12572_),
    .ZN(_12693_));
 AOI221_X2 _23127_ (.A(_12684_),
    .B1(_12690_),
    .B2(_12691_),
    .C1(_12692_),
    .C2(_12693_),
    .ZN(_12694_));
 MUX2_X1 _23128_ (.A(_12432_),
    .B(_12452_),
    .S(_12555_),
    .Z(_12695_));
 NAND2_X1 _23129_ (.A1(_12550_),
    .A2(_12695_),
    .ZN(_12696_));
 OAI21_X1 _23130_ (.A(_12558_),
    .B1(_12461_),
    .B2(_12494_),
    .ZN(_12697_));
 OAI22_X2 _23131_ (.A1(_12558_),
    .A2(_12599_),
    .B1(_12697_),
    .B2(_12614_),
    .ZN(_12698_));
 OAI221_X2 _23132_ (.A(_12696_),
    .B1(_12698_),
    .B2(_12619_),
    .C1(_12593_),
    .C2(_12536_),
    .ZN(_12699_));
 AOI21_X2 _23133_ (.A(_12699_),
    .B1(_12584_),
    .B2(_12557_),
    .ZN(_12700_));
 NOR2_X1 _23134_ (.A1(_12619_),
    .A2(_12616_),
    .ZN(_12701_));
 MUX2_X1 _23135_ (.A(_12439_),
    .B(_12412_),
    .S(_12555_),
    .Z(_12702_));
 AOI221_X2 _23136_ (.A(_12701_),
    .B1(_12702_),
    .B2(_12550_),
    .C1(_12557_),
    .C2(_12677_),
    .ZN(_12703_));
 NOR3_X2 _23137_ (.A1(_12694_),
    .A2(_12700_),
    .A3(_12703_),
    .ZN(_12704_));
 NAND3_X1 _23138_ (.A1(_12572_),
    .A2(_12631_),
    .A3(_12640_),
    .ZN(_12705_));
 NAND2_X1 _23139_ (.A1(_12488_),
    .A2(_12573_),
    .ZN(_12706_));
 AOI221_X2 _23140_ (.A(_12558_),
    .B1(_12452_),
    .B2(_12573_),
    .C1(_12706_),
    .C2(_12432_),
    .ZN(_12707_));
 NOR3_X1 _23141_ (.A1(_12572_),
    .A2(_12547_),
    .A3(_12707_),
    .ZN(_12708_));
 MUX2_X1 _23142_ (.A(_12439_),
    .B(_12412_),
    .S(_21229_),
    .Z(_12709_));
 OAI21_X1 _23143_ (.A(_12708_),
    .B1(_12709_),
    .B2(_12561_),
    .ZN(_12710_));
 MUX2_X1 _23144_ (.A(_12488_),
    .B(_12432_),
    .S(_12555_),
    .Z(_12711_));
 NAND2_X1 _23145_ (.A1(_12550_),
    .A2(_12711_),
    .ZN(_12712_));
 OAI221_X1 _23146_ (.A(_21234_),
    .B1(_12503_),
    .B2(_12504_),
    .C1(_12462_),
    .C2(_12499_),
    .ZN(_12713_));
 OAI21_X1 _23147_ (.A(_12713_),
    .B1(_12505_),
    .B2(_21234_),
    .ZN(_12714_));
 NAND4_X1 _23148_ (.A1(_12644_),
    .A2(_12591_),
    .A3(_12565_),
    .A4(_12714_),
    .ZN(_12715_));
 NAND4_X2 _23149_ (.A1(_12705_),
    .A2(_12710_),
    .A3(_12712_),
    .A4(_12715_),
    .ZN(_12716_));
 NAND2_X2 _23150_ (.A1(_12704_),
    .A2(_12716_),
    .ZN(_12717_));
 NOR4_X4 _23151_ (.A1(_12652_),
    .A2(_12670_),
    .A3(_12680_),
    .A4(_12717_),
    .ZN(_12718_));
 OAI21_X1 _23152_ (.A(_12609_),
    .B1(_12612_),
    .B2(_12718_),
    .ZN(_12719_));
 INV_X1 _23153_ (.A(_21239_),
    .ZN(_12720_));
 NOR3_X1 _23154_ (.A1(_12720_),
    .A2(_12161_),
    .A3(_12603_),
    .ZN(_12721_));
 AOI21_X2 _23155_ (.A(_12719_),
    .B1(_12721_),
    .B2(_12718_),
    .ZN(_12722_));
 AOI21_X2 _23156_ (.A(_12569_),
    .B1(_12161_),
    .B2(\g_reduce0[12].adder.a[0] ),
    .ZN(_12723_));
 AOI22_X4 _23157_ (.A1(_12198_),
    .A2(_12569_),
    .B1(_12722_),
    .B2(_12723_),
    .ZN(_00032_));
 NAND2_X4 _23158_ (.A1(_12157_),
    .A2(_12161_),
    .ZN(_12724_));
 INV_X1 _23159_ (.A(_12724_),
    .ZN(_12725_));
 AOI22_X4 _23160_ (.A1(\g_reduce0[12].adder.b[1] ),
    .A2(_12569_),
    .B1(_12725_),
    .B2(\g_reduce0[12].adder.a[1] ),
    .ZN(_12726_));
 INV_X1 _23161_ (.A(_21238_),
    .ZN(_12727_));
 MUX2_X1 _23162_ (.A(_12503_),
    .B(_12504_),
    .S(_12549_),
    .Z(_12728_));
 NAND2_X1 _23163_ (.A1(_12550_),
    .A2(_12728_),
    .ZN(_12729_));
 OAI21_X1 _23164_ (.A(_12729_),
    .B1(_12619_),
    .B2(_12604_),
    .ZN(_12730_));
 AOI21_X2 _23165_ (.A(_12730_),
    .B1(_12629_),
    .B2(_12557_),
    .ZN(_12731_));
 XNOR2_X1 _23166_ (.A(_12727_),
    .B(_12731_),
    .ZN(_12732_));
 OR4_X2 _23167_ (.A1(_12652_),
    .A2(_12670_),
    .A3(_12680_),
    .A4(_12717_),
    .ZN(_12733_));
 INV_X1 _23168_ (.A(_12603_),
    .ZN(_12734_));
 XNOR2_X1 _23169_ (.A(_12733_),
    .B(_12734_),
    .ZN(_12735_));
 INV_X2 _23170_ (.A(_12735_),
    .ZN(_21242_));
 MUX2_X1 _23171_ (.A(_12720_),
    .B(_12732_),
    .S(_21242_),
    .Z(_12736_));
 NAND2_X4 _23172_ (.A1(_12157_),
    .A2(_12611_),
    .ZN(_12737_));
 OAI21_X2 _23173_ (.A(_12726_),
    .B1(_12736_),
    .B2(_12737_),
    .ZN(_00039_));
 OAI22_X4 _23174_ (.A1(\g_reduce0[12].adder.b[2] ),
    .A2(_12157_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[2] ),
    .ZN(_12738_));
 OR2_X1 _23175_ (.A1(_12603_),
    .A2(_12732_),
    .ZN(_12739_));
 NOR2_X1 _23176_ (.A1(_12718_),
    .A2(_12739_),
    .ZN(_12740_));
 NOR2_X1 _23177_ (.A1(_12737_),
    .A2(_12740_),
    .ZN(_12741_));
 NOR2_X1 _23178_ (.A1(_12733_),
    .A2(_12732_),
    .ZN(_12742_));
 NAND2_X1 _23179_ (.A1(_12635_),
    .A2(_12651_),
    .ZN(_12743_));
 XNOR2_X1 _23180_ (.A(_12647_),
    .B(_12743_),
    .ZN(_12744_));
 OAI21_X1 _23181_ (.A(_12603_),
    .B1(_12742_),
    .B2(_12744_),
    .ZN(_12745_));
 AOI21_X2 _23182_ (.A(_12738_),
    .B1(_12741_),
    .B2(_12745_),
    .ZN(_00040_));
 NAND2_X1 _23183_ (.A1(\g_reduce0[12].adder.b[3] ),
    .A2(_12569_),
    .ZN(_12746_));
 BUF_X4 _23184_ (.A(_12157_),
    .Z(_12747_));
 OAI21_X1 _23185_ (.A(_12747_),
    .B1(_12611_),
    .B2(\g_reduce0[12].adder.a[3] ),
    .ZN(_12748_));
 NOR2_X2 _23186_ (.A1(_12727_),
    .A2(_12731_),
    .ZN(_12749_));
 NAND2_X1 _23187_ (.A1(_12647_),
    .A2(_12749_),
    .ZN(_12750_));
 XOR2_X1 _23188_ (.A(_12645_),
    .B(_12750_),
    .Z(_12751_));
 NOR3_X1 _23189_ (.A1(_12718_),
    .A2(_12734_),
    .A3(_12751_),
    .ZN(_12752_));
 AND2_X1 _23190_ (.A1(_12734_),
    .A2(_12744_),
    .ZN(_12753_));
 OAI21_X1 _23191_ (.A(_12611_),
    .B1(_12733_),
    .B2(_12739_),
    .ZN(_12754_));
 NOR3_X1 _23192_ (.A1(_12752_),
    .A2(_12753_),
    .A3(_12754_),
    .ZN(_12755_));
 OAI21_X2 _23193_ (.A(_12746_),
    .B1(_12748_),
    .B2(_12755_),
    .ZN(_00041_));
 INV_X1 _23194_ (.A(_12703_),
    .ZN(_12756_));
 XNOR2_X1 _23195_ (.A(_12652_),
    .B(_12756_),
    .ZN(_12757_));
 NOR2_X1 _23196_ (.A1(_12737_),
    .A2(_12757_),
    .ZN(_12758_));
 NOR2_X1 _23197_ (.A1(_12569_),
    .A2(_12161_),
    .ZN(_12759_));
 AND2_X1 _23198_ (.A1(_12759_),
    .A2(_12751_),
    .ZN(_12760_));
 MUX2_X1 _23199_ (.A(_12758_),
    .B(_12760_),
    .S(_12735_),
    .Z(_12761_));
 OAI22_X2 _23200_ (.A1(\g_reduce0[12].adder.b[4] ),
    .A2(_12747_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[4] ),
    .ZN(_12762_));
 NOR2_X1 _23201_ (.A1(_12761_),
    .A2(_12762_),
    .ZN(_00042_));
 OAI22_X4 _23202_ (.A1(\g_reduce0[12].adder.b[5] ),
    .A2(_12747_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[5] ),
    .ZN(_12763_));
 NAND4_X1 _23203_ (.A1(_12645_),
    .A2(_12647_),
    .A3(_12756_),
    .A4(_12749_),
    .ZN(_12764_));
 XOR2_X1 _23204_ (.A(_12694_),
    .B(_12764_),
    .Z(_12765_));
 NOR2_X1 _23205_ (.A1(_12737_),
    .A2(_12765_),
    .ZN(_12766_));
 MUX2_X1 _23206_ (.A(_12758_),
    .B(_12766_),
    .S(_21242_),
    .Z(_12767_));
 NOR2_X2 _23207_ (.A1(_12763_),
    .A2(_12767_),
    .ZN(_00043_));
 OAI22_X4 _23208_ (.A1(\g_reduce0[12].adder.b[6] ),
    .A2(_12747_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[6] ),
    .ZN(_12768_));
 AND2_X1 _23209_ (.A1(_12735_),
    .A2(_12766_),
    .ZN(_12769_));
 NOR3_X1 _23210_ (.A1(_12652_),
    .A2(_12694_),
    .A3(_12703_),
    .ZN(_12770_));
 XNOR2_X1 _23211_ (.A(_12700_),
    .B(_12770_),
    .ZN(_12771_));
 NOR3_X1 _23212_ (.A1(_12735_),
    .A2(_12737_),
    .A3(_12771_),
    .ZN(_12772_));
 NOR3_X1 _23213_ (.A1(_12768_),
    .A2(_12769_),
    .A3(_12772_),
    .ZN(_00044_));
 OAI22_X4 _23214_ (.A1(\g_reduce0[12].adder.b[7] ),
    .A2(_12747_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[7] ),
    .ZN(_12773_));
 NOR3_X1 _23215_ (.A1(_21242_),
    .A2(_12737_),
    .A3(_12771_),
    .ZN(_12774_));
 NAND4_X1 _23216_ (.A1(_12645_),
    .A2(_12647_),
    .A3(_12704_),
    .A4(_12749_),
    .ZN(_12775_));
 XOR2_X1 _23217_ (.A(_12716_),
    .B(_12775_),
    .Z(_12776_));
 NAND2_X1 _23218_ (.A1(_12759_),
    .A2(_12776_),
    .ZN(_12777_));
 NOR2_X1 _23219_ (.A1(_12735_),
    .A2(_12777_),
    .ZN(_12778_));
 NOR3_X1 _23220_ (.A1(_12773_),
    .A2(_12774_),
    .A3(_12778_),
    .ZN(_00045_));
 OAI22_X4 _23221_ (.A1(\g_reduce0[12].adder.b[8] ),
    .A2(_12747_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[8] ),
    .ZN(_12779_));
 NOR2_X1 _23222_ (.A1(_21242_),
    .A2(_12777_),
    .ZN(_12780_));
 NOR2_X1 _23223_ (.A1(_12652_),
    .A2(_12717_),
    .ZN(_12781_));
 XNOR2_X1 _23224_ (.A(_12680_),
    .B(_12781_),
    .ZN(_12782_));
 NOR3_X1 _23225_ (.A1(_12735_),
    .A2(_12737_),
    .A3(_12782_),
    .ZN(_12783_));
 NOR3_X1 _23226_ (.A1(_12779_),
    .A2(_12780_),
    .A3(_12783_),
    .ZN(_00046_));
 OAI22_X4 _23227_ (.A1(\g_reduce0[12].adder.b[9] ),
    .A2(_12157_),
    .B1(_12724_),
    .B2(\g_reduce0[12].adder.a[9] ),
    .ZN(_12784_));
 NOR3_X1 _23228_ (.A1(_21242_),
    .A2(_12737_),
    .A3(_12782_),
    .ZN(_12785_));
 NAND3_X1 _23229_ (.A1(_12645_),
    .A2(_12647_),
    .A3(_12749_),
    .ZN(_12786_));
 NOR3_X1 _23230_ (.A1(_12680_),
    .A2(_12717_),
    .A3(_12786_),
    .ZN(_12787_));
 XNOR2_X1 _23231_ (.A(_12670_),
    .B(_12787_),
    .ZN(_12788_));
 NOR3_X1 _23232_ (.A1(_12735_),
    .A2(_12737_),
    .A3(_12788_),
    .ZN(_12789_));
 NOR3_X1 _23233_ (.A1(_12784_),
    .A2(_12785_),
    .A3(_12789_),
    .ZN(_00047_));
 INV_X1 _23234_ (.A(_21246_),
    .ZN(_21240_));
 MUX2_X1 _23235_ (.A(\g_reduce0[12].adder.a[10] ),
    .B(_21245_),
    .S(_12611_),
    .Z(_12790_));
 MUX2_X2 _23236_ (.A(\g_reduce0[12].adder.b[10] ),
    .B(_12790_),
    .S(_12747_),
    .Z(_00033_));
 MUX2_X1 _23237_ (.A(\g_reduce0[12].adder.a[11] ),
    .B(_21253_),
    .S(_12611_),
    .Z(_12791_));
 MUX2_X2 _23238_ (.A(\g_reduce0[12].adder.b[11] ),
    .B(_12791_),
    .S(_12747_),
    .Z(_00034_));
 MUX2_X2 _23239_ (.A(_21121_),
    .B(_00486_),
    .S(_12205_),
    .Z(_12792_));
 NAND2_X1 _23240_ (.A1(_12549_),
    .A2(_21247_),
    .ZN(_12793_));
 XOR2_X1 _23241_ (.A(_12792_),
    .B(_12793_),
    .Z(_12794_));
 XOR2_X1 _23242_ (.A(_14070_),
    .B(_21257_),
    .Z(_12795_));
 MUX2_X1 _23243_ (.A(_12794_),
    .B(_12795_),
    .S(_12644_),
    .Z(_12796_));
 XOR2_X1 _23244_ (.A(_21252_),
    .B(_12796_),
    .Z(_12797_));
 MUX2_X1 _23245_ (.A(_12154_),
    .B(_12797_),
    .S(_12611_),
    .Z(_12798_));
 MUX2_X2 _23246_ (.A(_12158_),
    .B(_12798_),
    .S(_12747_),
    .Z(_00035_));
 INV_X1 _23247_ (.A(_14072_),
    .ZN(_14069_));
 MUX2_X1 _23248_ (.A(_21118_),
    .B(_00489_),
    .S(_12205_),
    .Z(_12799_));
 MUX2_X1 _23249_ (.A(_21124_),
    .B(_00481_),
    .S(_12205_),
    .Z(_12800_));
 NOR4_X1 _23250_ (.A1(_12555_),
    .A2(_21240_),
    .A3(_12792_),
    .A4(_12800_),
    .ZN(_12801_));
 XNOR2_X1 _23251_ (.A(_12799_),
    .B(_12801_),
    .ZN(_12802_));
 INV_X1 _23252_ (.A(_21249_),
    .ZN(_12803_));
 INV_X1 _23253_ (.A(_21250_),
    .ZN(_12804_));
 OAI21_X1 _23254_ (.A(_12803_),
    .B1(_12804_),
    .B2(_14072_),
    .ZN(_12805_));
 AOI21_X1 _23255_ (.A(_21256_),
    .B1(_12805_),
    .B2(_21257_),
    .ZN(_12806_));
 XNOR2_X1 _23256_ (.A(_21261_),
    .B(_12806_),
    .ZN(_12807_));
 MUX2_X1 _23257_ (.A(_12802_),
    .B(_12807_),
    .S(_12644_),
    .Z(_12808_));
 NAND2_X1 _23258_ (.A1(_12549_),
    .A2(_21248_),
    .ZN(_12809_));
 OAI21_X1 _23259_ (.A(_12809_),
    .B1(_12800_),
    .B2(_12549_),
    .ZN(_12810_));
 MUX2_X1 _23260_ (.A(_12810_),
    .B(_14071_),
    .S(_12644_),
    .Z(_21251_));
 NAND3_X1 _23261_ (.A1(_21244_),
    .A2(_12796_),
    .A3(_21251_),
    .ZN(_12811_));
 XNOR2_X1 _23262_ (.A(_12808_),
    .B(_12811_),
    .ZN(_12812_));
 MUX2_X1 _23263_ (.A(\g_reduce0[12].adder.a[13] ),
    .B(_12812_),
    .S(_12611_),
    .Z(_12813_));
 MUX2_X2 _23264_ (.A(\g_reduce0[12].adder.b[13] ),
    .B(_12813_),
    .S(_12747_),
    .Z(_00036_));
 OR2_X1 _23265_ (.A1(_12159_),
    .A2(_12193_),
    .ZN(_12814_));
 NAND2_X1 _23266_ (.A1(\g_reduce0[12].adder.a[14] ),
    .A2(_12814_),
    .ZN(_12815_));
 NOR3_X1 _23267_ (.A1(_12792_),
    .A2(_12793_),
    .A3(_12799_),
    .ZN(_12816_));
 AOI21_X1 _23268_ (.A(_21256_),
    .B1(_21257_),
    .B2(_14070_),
    .ZN(_12817_));
 INV_X1 _23269_ (.A(_12817_),
    .ZN(_12818_));
 AOI21_X1 _23270_ (.A(_21260_),
    .B1(_12818_),
    .B2(_21261_),
    .ZN(_12819_));
 MUX2_X1 _23271_ (.A(_12816_),
    .B(_12819_),
    .S(_12644_),
    .Z(_12820_));
 NAND3_X1 _23272_ (.A1(_21252_),
    .A2(_12796_),
    .A3(_12808_),
    .ZN(_12821_));
 XNOR2_X2 _23273_ (.A(_12820_),
    .B(_12821_),
    .ZN(_12822_));
 MUX2_X1 _23274_ (.A(_12814_),
    .B(_12815_),
    .S(_12822_),
    .Z(_12823_));
 OAI22_X1 _23275_ (.A1(_12159_),
    .A2(_12157_),
    .B1(_12161_),
    .B2(_12823_),
    .ZN(_12824_));
 NOR2_X1 _23276_ (.A1(\g_reduce0[12].adder.a[14] ),
    .A2(_12569_),
    .ZN(_12825_));
 NAND3_X1 _23277_ (.A1(_12159_),
    .A2(_12254_),
    .A3(_12822_),
    .ZN(_12826_));
 OR2_X1 _23278_ (.A1(_12254_),
    .A2(_12822_),
    .ZN(_12827_));
 NAND3_X1 _23279_ (.A1(_12611_),
    .A2(_12826_),
    .A3(_12827_),
    .ZN(_12828_));
 AOI21_X2 _23280_ (.A(_12824_),
    .B1(_12825_),
    .B2(_12828_),
    .ZN(_00037_));
 BUF_X2 _23281_ (.A(\g_reduce0[14].adder.a[11] ),
    .Z(_12829_));
 CLKBUF_X2 _23282_ (.A(\g_reduce0[14].adder.a[14] ),
    .Z(_12830_));
 OR2_X1 _23283_ (.A1(\g_reduce0[14].adder.a[10] ),
    .A2(\g_reduce0[14].adder.a[13] ),
    .ZN(_12831_));
 OR4_X1 _23284_ (.A1(_12829_),
    .A2(\g_reduce0[14].adder.a[12] ),
    .A3(_12830_),
    .A4(_12831_),
    .ZN(_12832_));
 CLKBUF_X3 _23285_ (.A(_12832_),
    .Z(_12833_));
 OR3_X1 _23286_ (.A1(\g_reduce0[14].adder.b[11] ),
    .A2(\g_reduce0[14].adder.b[10] ),
    .A3(\g_reduce0[14].adder.b[13] ),
    .ZN(_12834_));
 NOR3_X2 _23287_ (.A1(\g_reduce0[14].adder.b[12] ),
    .A2(\g_reduce0[14].adder.b[14] ),
    .A3(_12834_),
    .ZN(_12835_));
 CLKBUF_X3 _23288_ (.A(_12835_),
    .Z(_12836_));
 INV_X1 _23289_ (.A(_21308_),
    .ZN(_12837_));
 BUF_X4 _23290_ (.A(_21264_),
    .Z(_12838_));
 AOI21_X2 _23291_ (.A(_21263_),
    .B1(_21266_),
    .B2(_12838_),
    .ZN(_12839_));
 BUF_X2 _23292_ (.A(_21309_),
    .Z(_12840_));
 INV_X2 _23293_ (.A(_12840_),
    .ZN(_12841_));
 OAI21_X2 _23294_ (.A(_12837_),
    .B1(_12839_),
    .B2(_12841_),
    .ZN(_12842_));
 BUF_X1 _23295_ (.A(_21267_),
    .Z(_12843_));
 NAND3_X4 _23296_ (.A1(_12840_),
    .A2(_12838_),
    .A3(_12843_),
    .ZN(_12844_));
 INV_X1 _23297_ (.A(_12844_),
    .ZN(_12845_));
 INV_X1 _23298_ (.A(_21269_),
    .ZN(_12846_));
 INV_X2 _23299_ (.A(_21270_),
    .ZN(_12847_));
 OAI21_X2 _23300_ (.A(_12846_),
    .B1(_21302_),
    .B2(_12847_),
    .ZN(_12848_));
 AOI21_X4 _23301_ (.A(_12842_),
    .B1(_12845_),
    .B2(_12848_),
    .ZN(_12849_));
 INV_X4 _23302_ (.A(_21303_),
    .ZN(_12850_));
 NOR3_X1 _23303_ (.A1(_12850_),
    .A2(_12847_),
    .A3(_12844_),
    .ZN(_12851_));
 NOR2_X2 _23304_ (.A1(_12849_),
    .A2(_12851_),
    .ZN(_12852_));
 AND4_X2 _23305_ (.A1(_21273_),
    .A2(_21276_),
    .A3(_21279_),
    .A4(_21282_),
    .ZN(_12853_));
 AND3_X1 _23306_ (.A1(_21285_),
    .A2(_21288_),
    .A3(_21291_),
    .ZN(_12854_));
 AND2_X1 _23307_ (.A1(_21297_),
    .A2(_21300_),
    .ZN(_12855_));
 NAND4_X4 _23308_ (.A1(_21294_),
    .A2(_12853_),
    .A3(_12854_),
    .A4(_12855_),
    .ZN(_12856_));
 NAND2_X2 _23309_ (.A1(_12851_),
    .A2(_12856_),
    .ZN(_12857_));
 AND3_X1 _23310_ (.A1(_21294_),
    .A2(_12853_),
    .A3(_12854_),
    .ZN(_12858_));
 INV_X1 _23311_ (.A(_21296_),
    .ZN(_12859_));
 INV_X1 _23312_ (.A(_21297_),
    .ZN(_12860_));
 OAI21_X1 _23313_ (.A(_12859_),
    .B1(_21299_),
    .B2(_12860_),
    .ZN(_12861_));
 INV_X1 _23314_ (.A(_21275_),
    .ZN(_12862_));
 AOI21_X1 _23315_ (.A(_21278_),
    .B1(_21279_),
    .B2(_21281_),
    .ZN(_12863_));
 INV_X1 _23316_ (.A(_21276_),
    .ZN(_12864_));
 OAI21_X1 _23317_ (.A(_12862_),
    .B1(_12863_),
    .B2(_12864_),
    .ZN(_12865_));
 AOI221_X2 _23318_ (.A(_21272_),
    .B1(_12858_),
    .B2(_12861_),
    .C1(_12865_),
    .C2(_21273_),
    .ZN(_12866_));
 INV_X1 _23319_ (.A(_21284_),
    .ZN(_12867_));
 NAND3_X1 _23320_ (.A1(_21285_),
    .A2(_21288_),
    .A3(_21291_),
    .ZN(_12868_));
 INV_X1 _23321_ (.A(_21293_),
    .ZN(_12869_));
 AOI21_X1 _23322_ (.A(_21287_),
    .B1(_21290_),
    .B2(_21288_),
    .ZN(_12870_));
 INV_X1 _23323_ (.A(_21285_),
    .ZN(_12871_));
 OAI221_X2 _23324_ (.A(_12867_),
    .B1(_12868_),
    .B2(_12869_),
    .C1(_12870_),
    .C2(_12871_),
    .ZN(_12872_));
 NAND2_X2 _23325_ (.A1(_12853_),
    .A2(_12872_),
    .ZN(_12873_));
 AOI21_X4 _23326_ (.A(_12857_),
    .B1(_12866_),
    .B2(_12873_),
    .ZN(_12874_));
 OR2_X1 _23327_ (.A1(_12852_),
    .A2(_12874_),
    .ZN(_12875_));
 BUF_X4 _23328_ (.A(_12875_),
    .Z(_12876_));
 CLKBUF_X3 _23329_ (.A(_12876_),
    .Z(_12877_));
 OAI21_X1 _23330_ (.A(_12833_),
    .B1(_12836_),
    .B2(_12877_),
    .ZN(_12878_));
 MUX2_X1 _23331_ (.A(\g_reduce0[14].adder.a[15] ),
    .B(\g_reduce0[14].adder.b[15] ),
    .S(_12878_),
    .Z(_00054_));
 MUX2_X2 _23332_ (.A(_00492_),
    .B(_21301_),
    .S(_12877_),
    .Z(_21387_));
 INV_X1 _23333_ (.A(_21302_),
    .ZN(_12879_));
 AOI21_X1 _23334_ (.A(_21269_),
    .B1(_12879_),
    .B2(_21270_),
    .ZN(_12880_));
 OAI221_X2 _23335_ (.A(_12837_),
    .B1(_12880_),
    .B2(_12844_),
    .C1(_12839_),
    .C2(_12841_),
    .ZN(_12881_));
 CLKBUF_X3 _23336_ (.A(_21303_),
    .Z(_12882_));
 NAND3_X2 _23337_ (.A1(_12882_),
    .A2(_21270_),
    .A3(_12845_),
    .ZN(_12883_));
 NOR2_X1 _23338_ (.A1(\g_reduce0[14].adder.b[12] ),
    .A2(_00500_),
    .ZN(_12884_));
 NAND3_X1 _23339_ (.A1(_12881_),
    .A2(_12883_),
    .A3(_12884_),
    .ZN(_12885_));
 NAND3_X1 _23340_ (.A1(_12851_),
    .A2(_12856_),
    .A3(_12884_),
    .ZN(_12886_));
 AND2_X2 _23341_ (.A1(_12866_),
    .A2(_12873_),
    .ZN(_12887_));
 NOR2_X1 _23342_ (.A1(\g_reduce0[14].adder.a[12] ),
    .A2(_21265_),
    .ZN(_12888_));
 OAI21_X1 _23343_ (.A(_12888_),
    .B1(_12851_),
    .B2(_12849_),
    .ZN(_12889_));
 OAI221_X2 _23344_ (.A(_12885_),
    .B1(_12886_),
    .B2(_12887_),
    .C1(_12874_),
    .C2(_12889_),
    .ZN(_12890_));
 NAND3_X1 _23345_ (.A1(_12840_),
    .A2(_12838_),
    .A3(_12890_),
    .ZN(_12891_));
 INV_X2 _23346_ (.A(_21305_),
    .ZN(_12892_));
 NOR2_X2 _23347_ (.A1(\g_reduce0[14].adder.b[11] ),
    .A2(_00495_),
    .ZN(_12893_));
 INV_X1 _23348_ (.A(_21300_),
    .ZN(_12894_));
 NAND3_X1 _23349_ (.A1(_21294_),
    .A2(_12853_),
    .A3(_12854_),
    .ZN(_12895_));
 AND2_X1 _23350_ (.A1(_21273_),
    .A2(_12865_),
    .ZN(_12896_));
 INV_X1 _23351_ (.A(_21272_),
    .ZN(_12897_));
 INV_X1 _23352_ (.A(_21299_),
    .ZN(_12898_));
 AOI21_X1 _23353_ (.A(_21296_),
    .B1(_12898_),
    .B2(_21297_),
    .ZN(_12899_));
 OAI21_X1 _23354_ (.A(_12897_),
    .B1(_12895_),
    .B2(_12899_),
    .ZN(_12900_));
 AND2_X1 _23355_ (.A1(_12853_),
    .A2(_12872_),
    .ZN(_12901_));
 OAI33_X1 _23356_ (.A1(_12860_),
    .A2(_12894_),
    .A3(_12895_),
    .B1(_12896_),
    .B2(_12900_),
    .B3(_12901_),
    .ZN(_12902_));
 OR2_X1 _23357_ (.A1(_12829_),
    .A2(_21268_),
    .ZN(_12903_));
 NOR2_X1 _23358_ (.A1(_12883_),
    .A2(_12903_),
    .ZN(_12904_));
 NOR2_X1 _23359_ (.A1(_12829_),
    .A2(_21268_),
    .ZN(_12905_));
 MUX2_X1 _23360_ (.A(_12905_),
    .B(_12893_),
    .S(_12881_),
    .Z(_12906_));
 AOI222_X2 _23361_ (.A1(_12874_),
    .A2(_12893_),
    .B1(_12902_),
    .B2(_12904_),
    .C1(_12906_),
    .C2(_12883_),
    .ZN(_12907_));
 NAND3_X1 _23362_ (.A1(_12841_),
    .A2(_12892_),
    .A3(_12907_),
    .ZN(_12908_));
 BUF_X2 _23363_ (.A(_12852_),
    .Z(_12909_));
 BUF_X2 _23364_ (.A(_12874_),
    .Z(_12910_));
 OR2_X1 _23365_ (.A1(\g_reduce0[14].adder.a[13] ),
    .A2(_21262_),
    .ZN(_12911_));
 OR3_X1 _23366_ (.A1(_12909_),
    .A2(_12910_),
    .A3(_12911_),
    .ZN(_12912_));
 NOR2_X1 _23367_ (.A1(\g_reduce0[14].adder.b[13] ),
    .A2(_00503_),
    .ZN(_12913_));
 OAI21_X2 _23368_ (.A(_12913_),
    .B1(_12874_),
    .B2(_12852_),
    .ZN(_12914_));
 OR2_X1 _23369_ (.A1(_12874_),
    .A2(_12889_),
    .ZN(_12915_));
 OAI21_X1 _23370_ (.A(_12884_),
    .B1(_12874_),
    .B2(_12852_),
    .ZN(_12916_));
 NAND4_X2 _23371_ (.A1(_12912_),
    .A2(_12914_),
    .A3(_12915_),
    .A4(_12916_),
    .ZN(_12917_));
 AND2_X1 _23372_ (.A1(_12902_),
    .A2(_12904_),
    .ZN(_12918_));
 INV_X1 _23373_ (.A(_12893_),
    .ZN(_12919_));
 MUX2_X1 _23374_ (.A(_12903_),
    .B(_12919_),
    .S(_12881_),
    .Z(_12920_));
 NAND3_X1 _23375_ (.A1(_12851_),
    .A2(_12856_),
    .A3(_12893_),
    .ZN(_12921_));
 OAI221_X2 _23376_ (.A(_12892_),
    .B1(_12851_),
    .B2(_12920_),
    .C1(_12921_),
    .C2(_12887_),
    .ZN(_12922_));
 NOR2_X1 _23377_ (.A1(_12918_),
    .A2(_12922_),
    .ZN(_12923_));
 OAI221_X2 _23378_ (.A(_12891_),
    .B1(_12908_),
    .B2(_12917_),
    .C1(_12844_),
    .C2(_12923_),
    .ZN(_12924_));
 INV_X1 _23379_ (.A(_12838_),
    .ZN(_12925_));
 NAND4_X1 _23380_ (.A1(_12841_),
    .A2(_12925_),
    .A3(_12912_),
    .A4(_12914_),
    .ZN(_12926_));
 INV_X2 _23381_ (.A(_12843_),
    .ZN(_12927_));
 NAND2_X1 _23382_ (.A1(_12841_),
    .A2(_12927_),
    .ZN(_12928_));
 AND2_X1 _23383_ (.A1(_12912_),
    .A2(_12914_),
    .ZN(_12929_));
 OAI221_X2 _23384_ (.A(_12926_),
    .B1(_12928_),
    .B2(_12917_),
    .C1(_12841_),
    .C2(_12929_),
    .ZN(_12930_));
 OR2_X1 _23385_ (.A1(_12924_),
    .A2(_12930_),
    .ZN(_12931_));
 INV_X1 _23386_ (.A(_21301_),
    .ZN(_12932_));
 NOR2_X2 _23387_ (.A1(_00492_),
    .A2(_12932_),
    .ZN(_12933_));
 AND3_X1 _23388_ (.A1(_12851_),
    .A2(_12856_),
    .A3(_12933_),
    .ZN(_12934_));
 NAND2_X1 _23389_ (.A1(_00492_),
    .A2(_12932_),
    .ZN(_12935_));
 AOI21_X2 _23390_ (.A(_12935_),
    .B1(_12883_),
    .B2(_12881_),
    .ZN(_12936_));
 MUX2_X1 _23391_ (.A(_12934_),
    .B(_12936_),
    .S(_12887_),
    .Z(_12937_));
 NAND3_X1 _23392_ (.A1(_12881_),
    .A2(_12883_),
    .A3(_12933_),
    .ZN(_12938_));
 AND2_X1 _23393_ (.A1(_00492_),
    .A2(_12932_),
    .ZN(_12939_));
 OAI21_X1 _23394_ (.A(_12939_),
    .B1(_12851_),
    .B2(_12849_),
    .ZN(_12940_));
 AND2_X1 _23395_ (.A1(_12851_),
    .A2(_12856_),
    .ZN(_12941_));
 OAI21_X1 _23396_ (.A(_12938_),
    .B1(_12940_),
    .B2(_12941_),
    .ZN(_12942_));
 NAND3_X1 _23397_ (.A1(_12838_),
    .A2(_12843_),
    .A3(_21270_),
    .ZN(_12943_));
 OAI33_X1 _23398_ (.A1(_12925_),
    .A2(_12927_),
    .A3(_12907_),
    .B1(_12937_),
    .B2(_12942_),
    .B3(_12943_),
    .ZN(_12944_));
 NOR2_X1 _23399_ (.A1(_12838_),
    .A2(_12843_),
    .ZN(_12945_));
 MUX2_X1 _23400_ (.A(_12945_),
    .B(_12838_),
    .S(_12890_),
    .Z(_12946_));
 AND3_X1 _23401_ (.A1(_12915_),
    .A2(_12916_),
    .A3(_12907_),
    .ZN(_12947_));
 AOI22_X2 _23402_ (.A1(_12887_),
    .A2(_12936_),
    .B1(_12933_),
    .B2(_12910_),
    .ZN(_12948_));
 AOI221_X2 _23403_ (.A(_12847_),
    .B1(_12857_),
    .B2(_12936_),
    .C1(_12933_),
    .C2(_12852_),
    .ZN(_12949_));
 AOI21_X2 _23404_ (.A(_12838_),
    .B1(_12948_),
    .B2(_12949_),
    .ZN(_12950_));
 AOI211_X2 _23405_ (.A(_12944_),
    .B(_12946_),
    .C1(_12947_),
    .C2(_12950_),
    .ZN(_12951_));
 CLKBUF_X3 _23406_ (.A(_12951_),
    .Z(_12952_));
 BUF_X1 _23407_ (.A(_21306_),
    .Z(_12953_));
 INV_X1 _23408_ (.A(_12953_),
    .ZN(_12954_));
 CLKBUF_X3 _23409_ (.A(_12954_),
    .Z(_12955_));
 MUX2_X1 _23410_ (.A(_00498_),
    .B(_21277_),
    .S(_12876_),
    .Z(_12956_));
 NOR2_X1 _23411_ (.A1(_12955_),
    .A2(_12956_),
    .ZN(_12957_));
 OAI221_X2 _23412_ (.A(_00496_),
    .B1(_12849_),
    .B2(_12851_),
    .C1(_12857_),
    .C2(_12887_),
    .ZN(_12958_));
 OAI21_X1 _23413_ (.A(_21283_),
    .B1(_12909_),
    .B2(_12910_),
    .ZN(_12959_));
 AND2_X1 _23414_ (.A1(_12958_),
    .A2(_12959_),
    .ZN(_12960_));
 AOI21_X1 _23415_ (.A(_12957_),
    .B1(_12960_),
    .B2(_12955_),
    .ZN(_12961_));
 NAND2_X1 _23416_ (.A1(_12850_),
    .A2(_12961_),
    .ZN(_12962_));
 INV_X1 _23417_ (.A(_00499_),
    .ZN(_12963_));
 OR3_X1 _23418_ (.A1(_12963_),
    .A2(_12909_),
    .A3(_12874_),
    .ZN(_12964_));
 OAI21_X1 _23419_ (.A(_21280_),
    .B1(_12909_),
    .B2(_12910_),
    .ZN(_12965_));
 AND2_X1 _23420_ (.A1(_12964_),
    .A2(_12965_),
    .ZN(_12966_));
 INV_X1 _23421_ (.A(_00497_),
    .ZN(_12967_));
 OR3_X1 _23422_ (.A1(_12967_),
    .A2(_12909_),
    .A3(_12910_),
    .ZN(_12968_));
 OAI21_X1 _23423_ (.A(_21286_),
    .B1(_12909_),
    .B2(_12910_),
    .ZN(_12969_));
 AND2_X1 _23424_ (.A1(_12968_),
    .A2(_12969_),
    .ZN(_12970_));
 MUX2_X1 _23425_ (.A(_12966_),
    .B(_12970_),
    .S(_12955_),
    .Z(_12971_));
 OAI21_X1 _23426_ (.A(_12962_),
    .B1(_12971_),
    .B2(_12850_),
    .ZN(_12972_));
 MUX2_X1 _23427_ (.A(_00494_),
    .B(_21292_),
    .S(_12876_),
    .Z(_12973_));
 MUX2_X1 _23428_ (.A(_21298_),
    .B(_00491_),
    .S(_12876_),
    .Z(_12974_));
 MUX2_X1 _23429_ (.A(_12973_),
    .B(_12974_),
    .S(_12955_),
    .Z(_12975_));
 MUX2_X1 _23430_ (.A(_00490_),
    .B(_21295_),
    .S(_12876_),
    .Z(_12976_));
 NOR2_X1 _23431_ (.A1(_12953_),
    .A2(_12976_),
    .ZN(_12977_));
 INV_X1 _23432_ (.A(_00493_),
    .ZN(_12978_));
 OR3_X1 _23433_ (.A1(_12978_),
    .A2(_12909_),
    .A3(_12910_),
    .ZN(_12979_));
 OAI21_X1 _23434_ (.A(_21289_),
    .B1(_12909_),
    .B2(_12910_),
    .ZN(_12980_));
 AND2_X1 _23435_ (.A1(_12979_),
    .A2(_12980_),
    .ZN(_12981_));
 AOI21_X1 _23436_ (.A(_12977_),
    .B1(_12981_),
    .B2(_12953_),
    .ZN(_12982_));
 MUX2_X1 _23437_ (.A(_12975_),
    .B(_12982_),
    .S(_12850_),
    .Z(_12983_));
 OAI21_X1 _23438_ (.A(_12843_),
    .B1(_12918_),
    .B2(_12922_),
    .ZN(_12984_));
 NAND3_X1 _23439_ (.A1(_12892_),
    .A2(_12927_),
    .A3(_12907_),
    .ZN(_12985_));
 NAND2_X1 _23440_ (.A1(_12984_),
    .A2(_12985_),
    .ZN(_12986_));
 BUF_X4 _23441_ (.A(_12986_),
    .Z(_12987_));
 MUX2_X1 _23442_ (.A(_12972_),
    .B(_12983_),
    .S(_12987_),
    .Z(_12988_));
 NAND2_X1 _23443_ (.A1(_12850_),
    .A2(_12953_),
    .ZN(_12989_));
 INV_X1 _23444_ (.A(_00502_),
    .ZN(_12990_));
 INV_X1 _23445_ (.A(_21274_),
    .ZN(_12991_));
 MUX2_X1 _23446_ (.A(_12990_),
    .B(_12991_),
    .S(_12876_),
    .Z(_12992_));
 NAND2_X1 _23447_ (.A1(_12882_),
    .A2(_12992_),
    .ZN(_12993_));
 MUX2_X1 _23448_ (.A(_00501_),
    .B(_21271_),
    .S(_12876_),
    .Z(_12994_));
 OAI21_X1 _23449_ (.A(_12993_),
    .B1(_12994_),
    .B2(_12882_),
    .ZN(_12995_));
 OAI21_X1 _23450_ (.A(_12989_),
    .B1(_12995_),
    .B2(_12953_),
    .ZN(_12996_));
 NAND2_X1 _23451_ (.A1(_12952_),
    .A2(_12987_),
    .ZN(_12997_));
 OAI22_X1 _23452_ (.A1(_12952_),
    .A2(_12988_),
    .B1(_12996_),
    .B2(_12997_),
    .ZN(_12998_));
 NAND2_X1 _23453_ (.A1(_12931_),
    .A2(_12998_),
    .ZN(_21373_));
 INV_X1 _23454_ (.A(_21373_),
    .ZN(_21370_));
 NOR2_X1 _23455_ (.A1(_12850_),
    .A2(_12961_),
    .ZN(_12999_));
 MUX2_X1 _23456_ (.A(_12966_),
    .B(_12992_),
    .S(_12953_),
    .Z(_13000_));
 AOI21_X1 _23457_ (.A(_12999_),
    .B1(_13000_),
    .B2(_12850_),
    .ZN(_13001_));
 NAND2_X1 _23458_ (.A1(_12882_),
    .A2(_12982_),
    .ZN(_13002_));
 INV_X1 _23459_ (.A(_00494_),
    .ZN(_13003_));
 INV_X1 _23460_ (.A(_21292_),
    .ZN(_13004_));
 MUX2_X1 _23461_ (.A(_13003_),
    .B(_13004_),
    .S(_12876_),
    .Z(_13005_));
 MUX2_X1 _23462_ (.A(_12970_),
    .B(_13005_),
    .S(_12955_),
    .Z(_13006_));
 OAI21_X1 _23463_ (.A(_13002_),
    .B1(_13006_),
    .B2(_12882_),
    .ZN(_13007_));
 MUX2_X1 _23464_ (.A(_13001_),
    .B(_13007_),
    .S(_12987_),
    .Z(_13008_));
 NAND2_X1 _23465_ (.A1(_12882_),
    .A2(_12994_),
    .ZN(_13009_));
 NAND2_X1 _23466_ (.A1(_12955_),
    .A2(_13009_),
    .ZN(_13010_));
 OAI22_X1 _23467_ (.A1(_12952_),
    .A2(_13008_),
    .B1(_13010_),
    .B2(_12997_),
    .ZN(_13011_));
 NAND2_X1 _23468_ (.A1(_12931_),
    .A2(_13011_),
    .ZN(_14079_));
 INV_X1 _23469_ (.A(_14079_),
    .ZN(_14074_));
 INV_X1 _23470_ (.A(_12952_),
    .ZN(_13012_));
 AND2_X1 _23471_ (.A1(_12931_),
    .A2(_13012_),
    .ZN(_13013_));
 NAND2_X1 _23472_ (.A1(_12987_),
    .A2(_13013_),
    .ZN(_13014_));
 OR2_X1 _23473_ (.A1(_13010_),
    .A2(_13014_),
    .ZN(_21325_));
 INV_X1 _23474_ (.A(_21325_),
    .ZN(_21329_));
 OR2_X1 _23475_ (.A1(_12996_),
    .A2(_13014_),
    .ZN(_21318_));
 INV_X1 _23476_ (.A(_21318_),
    .ZN(_21322_));
 NOR2_X2 _23477_ (.A1(_12850_),
    .A2(_12953_),
    .ZN(_13015_));
 NAND2_X2 _23478_ (.A1(_12882_),
    .A2(_12953_),
    .ZN(_13016_));
 INV_X1 _23479_ (.A(_13016_),
    .ZN(_13017_));
 AOI22_X2 _23480_ (.A1(_12956_),
    .A2(_13015_),
    .B1(_13017_),
    .B2(_12994_),
    .ZN(_13018_));
 NAND2_X2 _23481_ (.A1(_12850_),
    .A2(_12954_),
    .ZN(_13019_));
 OR2_X1 _23482_ (.A1(_12992_),
    .A2(_13019_),
    .ZN(_13020_));
 NAND2_X1 _23483_ (.A1(_13018_),
    .A2(_13020_),
    .ZN(_13021_));
 OR2_X1 _23484_ (.A1(_13014_),
    .A2(_13021_),
    .ZN(_21353_));
 INV_X1 _23485_ (.A(_21353_),
    .ZN(_21357_));
 INV_X1 _23486_ (.A(_00498_),
    .ZN(_13022_));
 INV_X1 _23487_ (.A(_21277_),
    .ZN(_13023_));
 MUX2_X1 _23488_ (.A(_13022_),
    .B(_13023_),
    .S(_12877_),
    .Z(_13024_));
 MUX2_X1 _23489_ (.A(_13024_),
    .B(_12966_),
    .S(_12882_),
    .Z(_13025_));
 MUX2_X1 _23490_ (.A(_12995_),
    .B(_13025_),
    .S(_12955_),
    .Z(_13026_));
 MUX2_X1 _23491_ (.A(_13015_),
    .B(_13026_),
    .S(_12987_),
    .Z(_13027_));
 NAND2_X1 _23492_ (.A1(_13013_),
    .A2(_13027_),
    .ZN(_21332_));
 INV_X1 _23493_ (.A(_21332_),
    .ZN(_21336_));
 AOI21_X4 _23494_ (.A(_12927_),
    .B1(_12907_),
    .B2(_12892_),
    .ZN(_13028_));
 NOR3_X4 _23495_ (.A1(_12843_),
    .A2(_12918_),
    .A3(_12922_),
    .ZN(_13029_));
 NOR2_X2 _23496_ (.A1(_13028_),
    .A2(_13029_),
    .ZN(_13030_));
 NAND3_X1 _23497_ (.A1(_12955_),
    .A2(_13030_),
    .A3(_13009_),
    .ZN(_13031_));
 OAI21_X1 _23498_ (.A(_13031_),
    .B1(_13001_),
    .B2(_13030_),
    .ZN(_13032_));
 AND2_X1 _23499_ (.A1(_13013_),
    .A2(_13032_),
    .ZN(_21339_));
 INV_X1 _23500_ (.A(_21339_),
    .ZN(_21343_));
 OR2_X1 _23501_ (.A1(_13030_),
    .A2(_12972_),
    .ZN(_13033_));
 OAI21_X1 _23502_ (.A(_13033_),
    .B1(_12996_),
    .B2(_12987_),
    .ZN(_13034_));
 AND2_X1 _23503_ (.A1(_13013_),
    .A2(_13034_),
    .ZN(_21346_));
 INV_X1 _23504_ (.A(_21346_),
    .ZN(_21350_));
 AOI21_X2 _23505_ (.A(_13019_),
    .B1(_12969_),
    .B2(_12968_),
    .ZN(_13035_));
 NAND2_X1 _23506_ (.A1(_12882_),
    .A2(_12954_),
    .ZN(_13036_));
 AOI21_X2 _23507_ (.A(_13036_),
    .B1(_12980_),
    .B2(_12979_),
    .ZN(_13037_));
 AOI21_X2 _23508_ (.A(_12989_),
    .B1(_12965_),
    .B2(_12964_),
    .ZN(_13038_));
 AOI21_X2 _23509_ (.A(_13016_),
    .B1(_12959_),
    .B2(_12958_),
    .ZN(_13039_));
 OR4_X1 _23510_ (.A1(_13035_),
    .A2(_13037_),
    .A3(_13038_),
    .A4(_13039_),
    .ZN(_13040_));
 OR2_X1 _23511_ (.A1(_13030_),
    .A2(_13040_),
    .ZN(_13041_));
 OAI21_X1 _23512_ (.A(_13041_),
    .B1(_13021_),
    .B2(_12987_),
    .ZN(_13042_));
 AND2_X1 _23513_ (.A1(_13013_),
    .A2(_13042_),
    .ZN(_21363_));
 INV_X1 _23514_ (.A(_21363_),
    .ZN(_21367_));
 MUX2_X1 _23515_ (.A(_12960_),
    .B(_12981_),
    .S(_12955_),
    .Z(_13043_));
 MUX2_X1 _23516_ (.A(_13006_),
    .B(_13043_),
    .S(_12850_),
    .Z(_13044_));
 MUX2_X1 _23517_ (.A(_13026_),
    .B(_13044_),
    .S(_12987_),
    .Z(_13045_));
 NAND2_X1 _23518_ (.A1(_13012_),
    .A2(_13045_),
    .ZN(_13046_));
 OAI21_X2 _23519_ (.A(_13015_),
    .B1(_13029_),
    .B2(_13028_),
    .ZN(_13047_));
 OAI21_X1 _23520_ (.A(_13046_),
    .B1(_13047_),
    .B2(_13012_),
    .ZN(_13048_));
 NAND2_X1 _23521_ (.A1(_12931_),
    .A2(_13048_),
    .ZN(_21360_));
 INV_X1 _23522_ (.A(_21360_),
    .ZN(_21314_));
 BUF_X2 _23523_ (.A(_21327_),
    .Z(_13049_));
 XOR2_X2 _23524_ (.A(\g_reduce0[14].adder.b[15] ),
    .B(\g_reduce0[14].adder.a[15] ),
    .Z(_13050_));
 BUF_X4 _23525_ (.A(_13050_),
    .Z(_13051_));
 BUF_X4 _23526_ (.A(_13051_),
    .Z(_13052_));
 INV_X1 _23527_ (.A(_21320_),
    .ZN(_13053_));
 NAND2_X1 _23528_ (.A1(_13053_),
    .A2(_13051_),
    .ZN(_13054_));
 NOR3_X1 _23529_ (.A1(_13049_),
    .A2(_21355_),
    .A3(_13054_),
    .ZN(_13055_));
 CLKBUF_X3 _23530_ (.A(_21356_),
    .Z(_13056_));
 CLKBUF_X2 _23531_ (.A(_21335_),
    .Z(_13057_));
 INV_X1 _23532_ (.A(_13057_),
    .ZN(_13058_));
 INV_X1 _23533_ (.A(_21344_),
    .ZN(_13059_));
 BUF_X2 _23534_ (.A(_21342_),
    .Z(_13060_));
 AOI21_X1 _23535_ (.A(_13058_),
    .B1(_13059_),
    .B2(_13060_),
    .ZN(_13061_));
 OAI21_X1 _23536_ (.A(_13056_),
    .B1(_21334_),
    .B2(_13061_),
    .ZN(_13062_));
 OR3_X1 _23537_ (.A1(_21344_),
    .A2(_21334_),
    .A3(_21351_),
    .ZN(_13063_));
 INV_X1 _23538_ (.A(_21368_),
    .ZN(_13064_));
 AOI21_X1 _23539_ (.A(_21361_),
    .B1(_14080_),
    .B2(_21362_),
    .ZN(_13065_));
 BUF_X2 _23540_ (.A(_21366_),
    .Z(_13066_));
 OAI21_X1 _23541_ (.A(_13064_),
    .B1(_13065_),
    .B2(_13066_),
    .ZN(_13067_));
 BUF_X2 _23542_ (.A(_21349_),
    .Z(_13068_));
 INV_X2 _23543_ (.A(_13068_),
    .ZN(_13069_));
 AOI21_X1 _23544_ (.A(_13063_),
    .B1(_13067_),
    .B2(_13069_),
    .ZN(_13070_));
 OAI21_X1 _23545_ (.A(_13055_),
    .B1(_13062_),
    .B2(_13070_),
    .ZN(_13071_));
 BUF_X2 _23546_ (.A(_21321_),
    .Z(_13072_));
 INV_X1 _23547_ (.A(_13072_),
    .ZN(_13073_));
 NOR2_X1 _23548_ (.A1(_13049_),
    .A2(_21320_),
    .ZN(_13074_));
 NAND3_X1 _23549_ (.A1(_13073_),
    .A2(_13052_),
    .A3(_13074_),
    .ZN(_13075_));
 AND2_X1 _23550_ (.A1(_13071_),
    .A2(_13075_),
    .ZN(_13076_));
 BUF_X2 _23551_ (.A(_21328_),
    .Z(_13077_));
 INV_X2 _23552_ (.A(_13077_),
    .ZN(_13078_));
 MUX2_X1 _23553_ (.A(_21330_),
    .B(_13078_),
    .S(_13051_),
    .Z(_13079_));
 NOR2_X1 _23554_ (.A1(_13072_),
    .A2(_13077_),
    .ZN(_13080_));
 INV_X1 _23555_ (.A(_21358_),
    .ZN(_13081_));
 INV_X2 _23556_ (.A(_13056_),
    .ZN(_13082_));
 INV_X1 _23557_ (.A(_13060_),
    .ZN(_13083_));
 INV_X1 _23558_ (.A(_21341_),
    .ZN(_13084_));
 AOI21_X2 _23559_ (.A(_13057_),
    .B1(_13083_),
    .B2(_13084_),
    .ZN(_13085_));
 CLKBUF_X2 _23560_ (.A(_21337_),
    .Z(_13086_));
 OAI21_X1 _23561_ (.A(_13082_),
    .B1(_13085_),
    .B2(_13086_),
    .ZN(_13087_));
 BUF_X1 _23562_ (.A(_21348_),
    .Z(_13088_));
 OR3_X1 _23563_ (.A1(_13086_),
    .A2(_21341_),
    .A3(_13088_),
    .ZN(_13089_));
 INV_X1 _23564_ (.A(_21365_),
    .ZN(_13090_));
 AOI21_X1 _23565_ (.A(_21316_),
    .B1(_14076_),
    .B2(_21317_),
    .ZN(_13091_));
 INV_X1 _23566_ (.A(_13066_),
    .ZN(_13092_));
 OAI21_X2 _23567_ (.A(_13090_),
    .B1(_13091_),
    .B2(_13092_),
    .ZN(_13093_));
 AOI21_X1 _23568_ (.A(_13089_),
    .B1(_13093_),
    .B2(_13068_),
    .ZN(_13094_));
 OAI21_X2 _23569_ (.A(_13081_),
    .B1(_13087_),
    .B2(_13094_),
    .ZN(_13095_));
 AOI221_X1 _23570_ (.A(_13079_),
    .B1(_13080_),
    .B2(_13095_),
    .C1(_21323_),
    .C2(_13078_),
    .ZN(_13096_));
 AOI22_X1 _23571_ (.A1(_13049_),
    .A2(_13052_),
    .B1(_13076_),
    .B2(_13096_),
    .ZN(_13097_));
 OR2_X1 _23572_ (.A1(_21330_),
    .A2(_21323_),
    .ZN(_13098_));
 NOR2_X1 _23573_ (.A1(_13086_),
    .A2(_21341_),
    .ZN(_13099_));
 NOR2_X1 _23574_ (.A1(_13088_),
    .A2(_21365_),
    .ZN(_13100_));
 NAND2_X1 _23575_ (.A1(_13099_),
    .A2(_13100_),
    .ZN(_13101_));
 INV_X1 _23576_ (.A(_21316_),
    .ZN(_13102_));
 INV_X1 _23577_ (.A(_21317_),
    .ZN(_13103_));
 AOI21_X1 _23578_ (.A(_21310_),
    .B1(_14073_),
    .B2(_21311_),
    .ZN(_13104_));
 OAI21_X2 _23579_ (.A(_13102_),
    .B1(_13103_),
    .B2(_13104_),
    .ZN(_13105_));
 AOI21_X1 _23580_ (.A(_13101_),
    .B1(_13105_),
    .B2(_13066_),
    .ZN(_13106_));
 INV_X1 _23581_ (.A(_13099_),
    .ZN(_13107_));
 OR2_X1 _23582_ (.A1(_13068_),
    .A2(_13088_),
    .ZN(_13108_));
 OAI221_X2 _23583_ (.A(_13082_),
    .B1(_13107_),
    .B2(_13108_),
    .C1(_13085_),
    .C2(_13086_),
    .ZN(_13109_));
 OAI21_X1 _23584_ (.A(_13081_),
    .B1(_13106_),
    .B2(_13109_),
    .ZN(_13110_));
 AOI21_X2 _23585_ (.A(_13098_),
    .B1(_13110_),
    .B2(_13073_),
    .ZN(_13111_));
 XNOR2_X2 _23586_ (.A(\g_reduce0[14].adder.b[15] ),
    .B(\g_reduce0[14].adder.a[15] ),
    .ZN(_13112_));
 BUF_X4 _23587_ (.A(_13112_),
    .Z(_13113_));
 OAI21_X2 _23588_ (.A(_13113_),
    .B1(_13078_),
    .B2(_21330_),
    .ZN(_13114_));
 NOR2_X4 _23589_ (.A1(_13111_),
    .A2(_13114_),
    .ZN(_13115_));
 NOR2_X1 _23590_ (.A1(_13097_),
    .A2(_13115_),
    .ZN(_13116_));
 NAND2_X1 _23591_ (.A1(_13076_),
    .A2(_13096_),
    .ZN(_13117_));
 INV_X1 _23592_ (.A(_13049_),
    .ZN(_13118_));
 OAI21_X2 _23593_ (.A(_13117_),
    .B1(_13113_),
    .B2(_13118_),
    .ZN(_13119_));
 INV_X1 _23594_ (.A(_13074_),
    .ZN(_13120_));
 AOI21_X1 _23595_ (.A(_21355_),
    .B1(_21334_),
    .B2(_13056_),
    .ZN(_13121_));
 NOR2_X1 _23596_ (.A1(_21344_),
    .A2(_13083_),
    .ZN(_13122_));
 OR2_X1 _23597_ (.A1(_21344_),
    .A2(_21351_),
    .ZN(_13123_));
 AOI21_X1 _23598_ (.A(_13068_),
    .B1(_13066_),
    .B2(_13064_),
    .ZN(_13124_));
 NOR2_X1 _23599_ (.A1(_21361_),
    .A2(_21368_),
    .ZN(_13125_));
 AOI21_X1 _23600_ (.A(_21312_),
    .B1(_14078_),
    .B2(_21313_),
    .ZN(_13126_));
 INV_X1 _23601_ (.A(_21362_),
    .ZN(_13127_));
 OAI21_X1 _23602_ (.A(_13125_),
    .B1(_13126_),
    .B2(_13127_),
    .ZN(_13128_));
 AOI21_X2 _23603_ (.A(_13123_),
    .B1(_13124_),
    .B2(_13128_),
    .ZN(_13129_));
 NAND2_X1 _23604_ (.A1(_13057_),
    .A2(_13056_),
    .ZN(_13130_));
 OR3_X1 _23605_ (.A1(_13122_),
    .A2(_13129_),
    .A3(_13130_),
    .ZN(_13131_));
 AOI21_X1 _23606_ (.A(_13073_),
    .B1(_13121_),
    .B2(_13131_),
    .ZN(_13132_));
 OAI221_X2 _23607_ (.A(_13052_),
    .B1(_13120_),
    .B2(_13132_),
    .C1(_13049_),
    .C2(_13077_),
    .ZN(_13133_));
 NOR2_X1 _23608_ (.A1(_13119_),
    .A2(_13133_),
    .ZN(_13134_));
 AND2_X1 _23609_ (.A1(_12838_),
    .A2(_12890_),
    .ZN(_13135_));
 OAI221_X2 _23610_ (.A(_12914_),
    .B1(_12911_),
    .B2(_12876_),
    .C1(_12925_),
    .C2(_12927_),
    .ZN(_13136_));
 OAI21_X2 _23611_ (.A(_12840_),
    .B1(_13135_),
    .B2(_13136_),
    .ZN(_13137_));
 OR3_X2 _23612_ (.A1(_12840_),
    .A2(_13135_),
    .A3(_13136_),
    .ZN(_13138_));
 AOI211_X2 _23613_ (.A(_12951_),
    .B(_13047_),
    .C1(_13137_),
    .C2(_13138_),
    .ZN(_13139_));
 BUF_X4 _23614_ (.A(_13139_),
    .Z(_13140_));
 MUX2_X1 _23615_ (.A(_13116_),
    .B(_13134_),
    .S(_13140_),
    .Z(_13141_));
 BUF_X4 _23616_ (.A(_13141_),
    .Z(_13142_));
 NOR2_X1 _23617_ (.A1(_21355_),
    .A2(_13112_),
    .ZN(_13143_));
 OR2_X1 _23618_ (.A1(_13070_),
    .A2(_13062_),
    .ZN(_13144_));
 AOI22_X4 _23619_ (.A1(_13113_),
    .A2(_13095_),
    .B1(_13143_),
    .B2(_13144_),
    .ZN(_13145_));
 XNOR2_X2 _23620_ (.A(_13072_),
    .B(_13145_),
    .ZN(_13146_));
 NOR2_X1 _23621_ (.A1(_13112_),
    .A2(_13067_),
    .ZN(_13147_));
 AOI21_X4 _23622_ (.A(_13147_),
    .B1(_13093_),
    .B2(_13112_),
    .ZN(_13148_));
 XNOR2_X2 _23623_ (.A(_13069_),
    .B(_13148_),
    .ZN(_13149_));
 AOI21_X1 _23624_ (.A(_21351_),
    .B1(_13067_),
    .B2(_13069_),
    .ZN(_13150_));
 OAI21_X2 _23625_ (.A(_13059_),
    .B1(_13060_),
    .B2(_13150_),
    .ZN(_13151_));
 AOI21_X1 _23626_ (.A(_13088_),
    .B1(_13093_),
    .B2(_13068_),
    .ZN(_13152_));
 OR2_X1 _23627_ (.A1(_13083_),
    .A2(_13152_),
    .ZN(_13153_));
 NOR2_X1 _23628_ (.A1(_21341_),
    .A2(_13051_),
    .ZN(_13154_));
 AOI22_X4 _23629_ (.A1(_13051_),
    .A2(_13151_),
    .B1(_13153_),
    .B2(_13154_),
    .ZN(_13155_));
 XNOR2_X2 _23630_ (.A(_13058_),
    .B(_13155_),
    .ZN(_13156_));
 XOR2_X1 _23631_ (.A(_14076_),
    .B(_21317_),
    .Z(_13157_));
 XOR2_X1 _23632_ (.A(_14080_),
    .B(_21362_),
    .Z(_13158_));
 MUX2_X2 _23633_ (.A(_13157_),
    .B(_13158_),
    .S(_13051_),
    .Z(_13159_));
 MUX2_X2 _23634_ (.A(_21372_),
    .B(_21374_),
    .S(_13052_),
    .Z(_13160_));
 NOR2_X1 _23635_ (.A1(_13159_),
    .A2(_13160_),
    .ZN(_13161_));
 NAND4_X2 _23636_ (.A1(_13146_),
    .A2(_13149_),
    .A3(_13156_),
    .A4(_13161_),
    .ZN(_13162_));
 NOR2_X1 _23637_ (.A1(_13113_),
    .A2(_13162_),
    .ZN(_13163_));
 OAI21_X2 _23638_ (.A(_12952_),
    .B1(_12930_),
    .B2(_12924_),
    .ZN(_13164_));
 NAND3_X2 _23639_ (.A1(_12986_),
    .A2(_13018_),
    .A3(_13020_),
    .ZN(_13165_));
 AND2_X1 _23640_ (.A1(_12947_),
    .A2(_12950_),
    .ZN(_13166_));
 OR2_X1 _23641_ (.A1(_12944_),
    .A2(_12946_),
    .ZN(_13167_));
 OAI22_X4 _23642_ (.A1(_12924_),
    .A2(_12930_),
    .B1(_13166_),
    .B2(_13167_),
    .ZN(_13168_));
 OAI222_X2 _23643_ (.A1(_12973_),
    .A2(_12989_),
    .B1(_13016_),
    .B2(_12976_),
    .C1(_13019_),
    .C2(_12974_),
    .ZN(_13169_));
 NOR4_X2 _23644_ (.A1(_13028_),
    .A2(_13029_),
    .A3(_13038_),
    .A4(_13039_),
    .ZN(_13170_));
 NOR2_X2 _23645_ (.A1(_13035_),
    .A2(_13037_),
    .ZN(_13171_));
 AOI22_X4 _23646_ (.A1(_12987_),
    .A2(_13169_),
    .B1(_13170_),
    .B2(_13171_),
    .ZN(_13172_));
 OAI221_X2 _23647_ (.A(_13163_),
    .B1(_13164_),
    .B2(_13165_),
    .C1(_13168_),
    .C2(_13172_),
    .ZN(_13173_));
 NOR2_X1 _23648_ (.A1(_13052_),
    .A2(_13162_),
    .ZN(_13174_));
 AND4_X1 _23649_ (.A1(_12951_),
    .A2(_12986_),
    .A3(_13018_),
    .A4(_13020_),
    .ZN(_13175_));
 OR2_X1 _23650_ (.A1(_12976_),
    .A2(_13016_),
    .ZN(_13176_));
 NOR2_X1 _23651_ (.A1(_12882_),
    .A2(_12955_),
    .ZN(_13177_));
 INV_X1 _23652_ (.A(_13019_),
    .ZN(_13178_));
 OR3_X1 _23653_ (.A1(_21298_),
    .A2(_12909_),
    .A3(_12910_),
    .ZN(_13179_));
 NOR2_X2 _23654_ (.A1(_12909_),
    .A2(_12910_),
    .ZN(_13180_));
 OAI21_X1 _23655_ (.A(_13179_),
    .B1(_13180_),
    .B2(_00491_),
    .ZN(_13181_));
 AOI222_X2 _23656_ (.A1(_12984_),
    .A2(_12985_),
    .B1(_13005_),
    .B2(_13177_),
    .C1(_13178_),
    .C2(_13181_),
    .ZN(_13182_));
 AOI221_X2 _23657_ (.A(_12951_),
    .B1(_13030_),
    .B2(_13040_),
    .C1(_13176_),
    .C2(_13182_),
    .ZN(_13183_));
 OAI221_X2 _23658_ (.A(_13174_),
    .B1(_13175_),
    .B2(_13183_),
    .C1(_12924_),
    .C2(_12930_),
    .ZN(_13184_));
 NAND2_X1 _23659_ (.A1(_13051_),
    .A2(_13121_),
    .ZN(_13185_));
 NAND2_X1 _23660_ (.A1(_13053_),
    .A2(_13130_),
    .ZN(_13186_));
 OAI22_X2 _23661_ (.A1(_13072_),
    .A2(_13054_),
    .B1(_13185_),
    .B2(_13186_),
    .ZN(_13187_));
 NOR2_X1 _23662_ (.A1(_21358_),
    .A2(_21323_),
    .ZN(_13188_));
 OAI21_X1 _23663_ (.A(_13188_),
    .B1(_13109_),
    .B2(_13106_),
    .ZN(_13189_));
 INV_X1 _23664_ (.A(_21323_),
    .ZN(_13190_));
 AOI21_X1 _23665_ (.A(_13051_),
    .B1(_13190_),
    .B2(_13072_),
    .ZN(_13191_));
 NOR2_X1 _23666_ (.A1(_21320_),
    .A2(_13185_),
    .ZN(_13192_));
 OR2_X2 _23667_ (.A1(_13122_),
    .A2(_13129_),
    .ZN(_13193_));
 AOI221_X2 _23668_ (.A(_13187_),
    .B1(_13189_),
    .B2(_13191_),
    .C1(_13192_),
    .C2(_13193_),
    .ZN(_13194_));
 XNOR2_X2 _23669_ (.A(_13077_),
    .B(_13194_),
    .ZN(_13195_));
 NAND2_X1 _23670_ (.A1(_21334_),
    .A2(_13052_),
    .ZN(_13196_));
 NOR2_X1 _23671_ (.A1(_13051_),
    .A2(_13107_),
    .ZN(_13197_));
 NAND2_X1 _23672_ (.A1(_13060_),
    .A2(_13108_),
    .ZN(_13198_));
 INV_X1 _23673_ (.A(_13100_),
    .ZN(_13199_));
 AOI21_X1 _23674_ (.A(_13199_),
    .B1(_13105_),
    .B2(_13066_),
    .ZN(_13200_));
 OAI21_X2 _23675_ (.A(_13197_),
    .B1(_13198_),
    .B2(_13200_),
    .ZN(_13201_));
 NAND2_X2 _23676_ (.A1(_13196_),
    .A2(_13201_),
    .ZN(_13202_));
 AOI21_X2 _23677_ (.A(_13058_),
    .B1(_13086_),
    .B2(_13113_),
    .ZN(_13203_));
 INV_X1 _23678_ (.A(_13203_),
    .ZN(_13204_));
 AOI21_X4 _23679_ (.A(_13204_),
    .B1(_13193_),
    .B2(_13052_),
    .ZN(_13205_));
 OAI21_X4 _23680_ (.A(_13056_),
    .B1(_13202_),
    .B2(_13205_),
    .ZN(_13206_));
 AND2_X2 _23681_ (.A1(_13196_),
    .A2(_13201_),
    .ZN(_13207_));
 NOR2_X1 _23682_ (.A1(_13122_),
    .A2(_13129_),
    .ZN(_13208_));
 OAI21_X4 _23683_ (.A(_13203_),
    .B1(_13208_),
    .B2(_13113_),
    .ZN(_13209_));
 NAND3_X4 _23684_ (.A1(_13082_),
    .A2(_13207_),
    .A3(_13209_),
    .ZN(_13210_));
 NOR3_X1 _23685_ (.A1(_13069_),
    .A2(_13090_),
    .A3(_13051_),
    .ZN(_13211_));
 NOR3_X1 _23686_ (.A1(_13069_),
    .A2(_13092_),
    .A3(_13050_),
    .ZN(_13212_));
 AOI221_X2 _23687_ (.A(_13211_),
    .B1(_13212_),
    .B2(_13105_),
    .C1(_13088_),
    .C2(_13112_),
    .ZN(_13213_));
 OR2_X1 _23688_ (.A1(_21351_),
    .A2(_13112_),
    .ZN(_13214_));
 AND2_X1 _23689_ (.A1(_13128_),
    .A2(_13124_),
    .ZN(_13215_));
 OAI21_X2 _23690_ (.A(_13213_),
    .B1(_13214_),
    .B2(_13215_),
    .ZN(_13216_));
 XNOR2_X2 _23691_ (.A(_13060_),
    .B(_13216_),
    .ZN(_13217_));
 OR2_X1 _23692_ (.A1(_13127_),
    .A2(_13126_),
    .ZN(_13218_));
 NOR2_X1 _23693_ (.A1(_21361_),
    .A2(_13112_),
    .ZN(_13219_));
 AOI22_X2 _23694_ (.A1(_13112_),
    .A2(_13105_),
    .B1(_13218_),
    .B2(_13219_),
    .ZN(_13220_));
 XNOR2_X2 _23695_ (.A(_13066_),
    .B(_13220_),
    .ZN(_13221_));
 AND2_X1 _23696_ (.A1(_14077_),
    .A2(_13113_),
    .ZN(_13222_));
 AOI21_X4 _23697_ (.A(_13222_),
    .B1(_13052_),
    .B2(_14081_),
    .ZN(_13223_));
 INV_X1 _23698_ (.A(_13159_),
    .ZN(_13224_));
 AOI21_X1 _23699_ (.A(_13221_),
    .B1(_13223_),
    .B2(_13224_),
    .ZN(_13225_));
 XNOR2_X2 _23700_ (.A(_13068_),
    .B(_13148_),
    .ZN(_13226_));
 OAI21_X2 _23701_ (.A(_13217_),
    .B1(_13225_),
    .B2(_13226_),
    .ZN(_13227_));
 AOI22_X4 _23702_ (.A1(_13206_),
    .A2(_13210_),
    .B1(_13227_),
    .B2(_13156_),
    .ZN(_13228_));
 XNOR2_X2 _23703_ (.A(_13073_),
    .B(_13145_),
    .ZN(_13229_));
 OAI21_X4 _23704_ (.A(_13195_),
    .B1(_13228_),
    .B2(_13229_),
    .ZN(_13230_));
 AOI211_X2 _23705_ (.A(_13115_),
    .B(_13230_),
    .C1(_13133_),
    .C2(_13140_),
    .ZN(_13231_));
 AND3_X2 _23706_ (.A1(_13173_),
    .A2(_13184_),
    .A3(_13231_),
    .ZN(_13232_));
 NOR2_X4 _23707_ (.A1(_13142_),
    .A2(_13232_),
    .ZN(_21375_));
 INV_X2 _23708_ (.A(_21375_),
    .ZN(_21378_));
 CLKBUF_X2 _23709_ (.A(_21381_),
    .Z(_13233_));
 INV_X1 _23710_ (.A(_13233_),
    .ZN(_13234_));
 OR2_X1 _23711_ (.A1(_13111_),
    .A2(_13114_),
    .ZN(_13235_));
 NAND3_X1 _23712_ (.A1(_13234_),
    .A2(_13097_),
    .A3(_13235_),
    .ZN(_13236_));
 XNOR2_X2 _23713_ (.A(_13057_),
    .B(_13155_),
    .ZN(_13237_));
 NOR2_X1 _23714_ (.A1(_13159_),
    .A2(_13221_),
    .ZN(_13238_));
 AND3_X2 _23715_ (.A1(_13149_),
    .A2(_13217_),
    .A3(_13238_),
    .ZN(_13239_));
 AOI211_X2 _23716_ (.A(_13237_),
    .B(_13239_),
    .C1(_13210_),
    .C2(_13206_),
    .ZN(_13240_));
 XNOR2_X2 _23717_ (.A(_13078_),
    .B(_13194_),
    .ZN(_13241_));
 NOR2_X2 _23718_ (.A1(_13229_),
    .A2(_13241_),
    .ZN(_13242_));
 AOI21_X1 _23719_ (.A(_13236_),
    .B1(_13240_),
    .B2(_13242_),
    .ZN(_13243_));
 NAND2_X1 _23720_ (.A1(_13071_),
    .A2(_13075_),
    .ZN(_13244_));
 OR3_X1 _23721_ (.A1(_13233_),
    .A2(_13244_),
    .A3(_13133_),
    .ZN(_13245_));
 AOI211_X2 _23722_ (.A(_12952_),
    .B(_13245_),
    .C1(_13240_),
    .C2(_13242_),
    .ZN(_13246_));
 AOI21_X2 _23723_ (.A(_13047_),
    .B1(_13137_),
    .B2(_13138_),
    .ZN(_13247_));
 MUX2_X1 _23724_ (.A(_13243_),
    .B(_13246_),
    .S(_13247_),
    .Z(_13248_));
 AND3_X1 _23725_ (.A1(_13234_),
    .A2(_13097_),
    .A3(_13235_),
    .ZN(_13249_));
 NAND3_X1 _23726_ (.A1(_13149_),
    .A2(_13217_),
    .A3(_13238_),
    .ZN(_13250_));
 NOR3_X4 _23727_ (.A1(_13056_),
    .A2(_13202_),
    .A3(_13205_),
    .ZN(_13251_));
 AOI21_X4 _23728_ (.A(_13082_),
    .B1(_13207_),
    .B2(_13209_),
    .ZN(_13252_));
 OAI211_X2 _23729_ (.A(_13156_),
    .B(_13250_),
    .C1(_13251_),
    .C2(_13252_),
    .ZN(_13253_));
 NAND2_X2 _23730_ (.A1(_13146_),
    .A2(_13195_),
    .ZN(_13254_));
 OAI211_X2 _23731_ (.A(_12952_),
    .B(_13249_),
    .C1(_13253_),
    .C2(_13254_),
    .ZN(_13255_));
 NAND2_X1 _23732_ (.A1(_13097_),
    .A2(_13235_),
    .ZN(_13256_));
 NAND3_X1 _23733_ (.A1(_13233_),
    .A2(_12952_),
    .A3(_13256_),
    .ZN(_13257_));
 NAND2_X1 _23734_ (.A1(_13233_),
    .A2(_13256_),
    .ZN(_13258_));
 OAI211_X2 _23735_ (.A(_13255_),
    .B(_13257_),
    .C1(_13247_),
    .C2(_13258_),
    .ZN(_13259_));
 NAND2_X1 _23736_ (.A1(_13206_),
    .A2(_13210_),
    .ZN(_13260_));
 NAND3_X2 _23737_ (.A1(_13156_),
    .A2(_13260_),
    .A3(_13242_),
    .ZN(_13261_));
 OR2_X1 _23738_ (.A1(_13244_),
    .A2(_13133_),
    .ZN(_13262_));
 NAND2_X1 _23739_ (.A1(_13233_),
    .A2(_13262_),
    .ZN(_13263_));
 OAI21_X1 _23740_ (.A(_12841_),
    .B1(_13135_),
    .B2(_13136_),
    .ZN(_13264_));
 OR3_X1 _23741_ (.A1(_12841_),
    .A2(_13135_),
    .A3(_13136_),
    .ZN(_13265_));
 NAND4_X2 _23742_ (.A1(_12987_),
    .A2(_13015_),
    .A3(_13264_),
    .A4(_13265_),
    .ZN(_13266_));
 OAI33_X1 _23743_ (.A1(_13234_),
    .A2(_13239_),
    .A3(_13261_),
    .B1(_13263_),
    .B2(_13266_),
    .B3(_12952_),
    .ZN(_13267_));
 NOR3_X4 _23744_ (.A1(_13248_),
    .A2(_13259_),
    .A3(_13267_),
    .ZN(_00616_));
 INV_X2 _23745_ (.A(_00616_),
    .ZN(_21401_));
 INV_X1 _23746_ (.A(_13256_),
    .ZN(_00617_));
 INV_X1 _23747_ (.A(_13262_),
    .ZN(_00618_));
 MUX2_X1 _23748_ (.A(_00617_),
    .B(_00618_),
    .S(_13140_),
    .Z(_00619_));
 CLKBUF_X3 _23749_ (.A(_00619_),
    .Z(_00620_));
 BUF_X4 _23750_ (.A(_00620_),
    .Z(_00621_));
 CLKBUF_X2 _23751_ (.A(_21377_),
    .Z(_00622_));
 INV_X1 _23752_ (.A(_00622_),
    .ZN(_00623_));
 CLKBUF_X3 _23753_ (.A(_00623_),
    .Z(_00624_));
 AND2_X1 _23754_ (.A1(_21372_),
    .A2(_13113_),
    .ZN(_00625_));
 AOI21_X4 _23755_ (.A(_00625_),
    .B1(_13052_),
    .B2(_21374_),
    .ZN(_00626_));
 NOR2_X1 _23756_ (.A1(_00624_),
    .A2(_00626_),
    .ZN(_00627_));
 OAI221_X2 _23757_ (.A(_13113_),
    .B1(_13165_),
    .B2(_13164_),
    .C1(_13172_),
    .C2(_13168_),
    .ZN(_00628_));
 OAI221_X2 _23758_ (.A(_13052_),
    .B1(_13183_),
    .B2(_13175_),
    .C1(_12930_),
    .C2(_12924_),
    .ZN(_00629_));
 AND2_X1 _23759_ (.A1(_00628_),
    .A2(_00629_),
    .ZN(_00630_));
 AOI21_X1 _23760_ (.A(_00627_),
    .B1(_00630_),
    .B2(_00624_),
    .ZN(_00631_));
 MUX2_X2 _23761_ (.A(_13256_),
    .B(_13262_),
    .S(_13140_),
    .Z(_00632_));
 NOR2_X1 _23762_ (.A1(_13254_),
    .A2(_13253_),
    .ZN(_00633_));
 XNOR2_X1 _23763_ (.A(_13234_),
    .B(_00633_),
    .ZN(_00634_));
 NOR2_X2 _23764_ (.A1(_00632_),
    .A2(_00634_),
    .ZN(_00635_));
 NOR2_X4 _23765_ (.A1(_13252_),
    .A2(_13251_),
    .ZN(_00636_));
 NOR3_X4 _23766_ (.A1(_13237_),
    .A2(_00636_),
    .A3(_13254_),
    .ZN(_00637_));
 OR2_X2 _23767_ (.A1(_13229_),
    .A2(_13228_),
    .ZN(_00638_));
 AND3_X2 _23768_ (.A1(_13173_),
    .A2(_13184_),
    .A3(_00638_),
    .ZN(_00639_));
 OAI21_X1 _23769_ (.A(_13238_),
    .B1(_13223_),
    .B2(_13160_),
    .ZN(_00640_));
 AND3_X1 _23770_ (.A1(_13149_),
    .A2(_13217_),
    .A3(_00640_),
    .ZN(_00641_));
 NOR3_X1 _23771_ (.A1(_13237_),
    .A2(_00636_),
    .A3(_00641_),
    .ZN(_00642_));
 OR2_X2 _23772_ (.A1(_13254_),
    .A2(_00642_),
    .ZN(_00643_));
 AOI21_X4 _23773_ (.A(_13261_),
    .B1(_00620_),
    .B2(_00643_),
    .ZN(_00644_));
 AOI22_X4 _23774_ (.A1(_13239_),
    .A2(_00637_),
    .B1(_00639_),
    .B2(_00644_),
    .ZN(_00645_));
 NAND2_X2 _23775_ (.A1(_00635_),
    .A2(_00645_),
    .ZN(_00646_));
 BUF_X2 _23776_ (.A(_14083_),
    .Z(_00647_));
 INV_X1 _23777_ (.A(_00647_),
    .ZN(_00648_));
 CLKBUF_X3 _23778_ (.A(_00648_),
    .Z(_00649_));
 INV_X1 _23779_ (.A(_13133_),
    .ZN(_00650_));
 OR2_X1 _23780_ (.A1(_12952_),
    .A2(_00650_),
    .ZN(_00651_));
 OAI21_X1 _23781_ (.A(_13235_),
    .B1(_13266_),
    .B2(_00651_),
    .ZN(_00652_));
 CLKBUF_X3 _23782_ (.A(_00652_),
    .Z(_00653_));
 XNOR2_X2 _23783_ (.A(_13119_),
    .B(_13139_),
    .ZN(_00654_));
 AOI22_X4 _23784_ (.A1(_00628_),
    .A2(_00629_),
    .B1(_13230_),
    .B2(_00654_),
    .ZN(_00655_));
 OR3_X1 _23785_ (.A1(_00649_),
    .A2(_00653_),
    .A3(_00655_),
    .ZN(_00656_));
 OAI22_X2 _23786_ (.A1(_00621_),
    .A2(_00631_),
    .B1(_00646_),
    .B2(_00656_),
    .ZN(_00657_));
 CLKBUF_X3 _23787_ (.A(_00622_),
    .Z(_00658_));
 MUX2_X1 _23788_ (.A(_14081_),
    .B(_14077_),
    .S(_13113_),
    .Z(_00659_));
 BUF_X4 _23789_ (.A(_00632_),
    .Z(_00660_));
 NAND3_X1 _23790_ (.A1(_00658_),
    .A2(_00659_),
    .A3(_00660_),
    .ZN(_00661_));
 OAI21_X1 _23791_ (.A(_00660_),
    .B1(_13160_),
    .B2(_00658_),
    .ZN(_00662_));
 NAND3_X1 _23792_ (.A1(_13162_),
    .A2(_13195_),
    .A3(_00638_),
    .ZN(_00663_));
 AND4_X1 _23793_ (.A1(_00647_),
    .A2(_00630_),
    .A3(_00620_),
    .A4(_00663_),
    .ZN(_00664_));
 NAND2_X1 _23794_ (.A1(_00647_),
    .A2(_00626_),
    .ZN(_00665_));
 AOI21_X4 _23795_ (.A(_00664_),
    .B1(_00665_),
    .B2(_21378_),
    .ZN(_00666_));
 OAI21_X1 _23796_ (.A(_00662_),
    .B1(_00666_),
    .B2(_00646_),
    .ZN(_00667_));
 AND3_X1 _23797_ (.A1(_00657_),
    .A2(_00661_),
    .A3(_00667_),
    .ZN(_21383_));
 NOR4_X4 _23798_ (.A1(_12829_),
    .A2(\g_reduce0[14].adder.a[12] ),
    .A3(_12830_),
    .A4(_12831_),
    .ZN(_00668_));
 AND2_X1 _23799_ (.A1(_12832_),
    .A2(_12836_),
    .ZN(_00669_));
 AOI22_X1 _23800_ (.A1(\g_reduce0[14].adder.b[0] ),
    .A2(_00668_),
    .B1(_00669_),
    .B2(\g_reduce0[14].adder.a[0] ),
    .ZN(_00670_));
 INV_X1 _23801_ (.A(_21386_),
    .ZN(_00671_));
 INV_X1 _23802_ (.A(_21379_),
    .ZN(_00672_));
 CLKBUF_X3 _23803_ (.A(_00616_),
    .Z(_00673_));
 AOI21_X4 _23804_ (.A(_13115_),
    .B1(_13140_),
    .B2(_13133_),
    .ZN(_00674_));
 NAND2_X1 _23805_ (.A1(_13239_),
    .A2(_00637_),
    .ZN(_00675_));
 NAND2_X1 _23806_ (.A1(_00674_),
    .A2(_00675_),
    .ZN(_00676_));
 AOI21_X2 _23807_ (.A(_00676_),
    .B1(_00644_),
    .B2(_00639_),
    .ZN(_00677_));
 NOR2_X2 _23808_ (.A1(_13142_),
    .A2(_00677_),
    .ZN(_00678_));
 NOR3_X1 _23809_ (.A1(_00672_),
    .A2(_00673_),
    .A3(_00678_),
    .ZN(_00679_));
 OAI21_X1 _23810_ (.A(_00657_),
    .B1(_00679_),
    .B2(_00660_),
    .ZN(_00680_));
 NAND2_X1 _23811_ (.A1(_00661_),
    .A2(_00667_),
    .ZN(_00681_));
 MUX2_X1 _23812_ (.A(_00657_),
    .B(_00680_),
    .S(_00681_),
    .Z(_00682_));
 CLKBUF_X3 _23813_ (.A(_00621_),
    .Z(_00683_));
 AOI21_X2 _23814_ (.A(_00683_),
    .B1(_21375_),
    .B2(_00624_),
    .ZN(_00684_));
 NOR2_X1 _23815_ (.A1(_00653_),
    .A2(_00655_),
    .ZN(_00685_));
 NOR3_X1 _23816_ (.A1(_13224_),
    .A2(_00638_),
    .A3(_00632_),
    .ZN(_00686_));
 XNOR2_X2 _23817_ (.A(_13097_),
    .B(_13140_),
    .ZN(_00687_));
 NOR4_X1 _23818_ (.A1(_00653_),
    .A2(_00687_),
    .A3(_13224_),
    .A4(_13195_),
    .ZN(_00688_));
 INV_X1 _23819_ (.A(_13221_),
    .ZN(_00689_));
 NOR3_X1 _23820_ (.A1(_13229_),
    .A2(_13226_),
    .A3(_13237_),
    .ZN(_00690_));
 XNOR2_X1 _23821_ (.A(_13083_),
    .B(_13216_),
    .ZN(_00691_));
 AOI22_X2 _23822_ (.A1(_13206_),
    .A2(_13210_),
    .B1(_00691_),
    .B2(_13156_),
    .ZN(_00692_));
 OAI21_X2 _23823_ (.A(_13195_),
    .B1(_00692_),
    .B2(_13229_),
    .ZN(_00693_));
 OR2_X1 _23824_ (.A1(_00690_),
    .A2(_00693_),
    .ZN(_00694_));
 AOI211_X2 _23825_ (.A(_00652_),
    .B(_00689_),
    .C1(_00694_),
    .C2(_00654_),
    .ZN(_00695_));
 OR3_X1 _23826_ (.A1(_00686_),
    .A2(_00688_),
    .A3(_00695_),
    .ZN(_00696_));
 MUX2_X1 _23827_ (.A(_00685_),
    .B(_00696_),
    .S(_21401_),
    .Z(_00697_));
 NOR2_X1 _23828_ (.A1(_00649_),
    .A2(_00697_),
    .ZN(_00698_));
 CLKBUF_X3 _23829_ (.A(_00647_),
    .Z(_00699_));
 NOR2_X1 _23830_ (.A1(_00626_),
    .A2(_13195_),
    .ZN(_00700_));
 MUX2_X1 _23831_ (.A(_13223_),
    .B(_00700_),
    .S(_13119_),
    .Z(_00701_));
 AND3_X1 _23832_ (.A1(_13140_),
    .A2(_00650_),
    .A3(_00701_),
    .ZN(_00702_));
 MUX2_X1 _23833_ (.A(_13223_),
    .B(_00700_),
    .S(_13097_),
    .Z(_00703_));
 NOR2_X1 _23834_ (.A1(_13115_),
    .A2(_13140_),
    .ZN(_00704_));
 NOR2_X1 _23835_ (.A1(_00626_),
    .A2(_00638_),
    .ZN(_00705_));
 AOI221_X2 _23836_ (.A(_00702_),
    .B1(_00703_),
    .B2(_00704_),
    .C1(_00705_),
    .C2(_00620_),
    .ZN(_00706_));
 NAND2_X1 _23837_ (.A1(_13223_),
    .A2(_13231_),
    .ZN(_00707_));
 NAND2_X1 _23838_ (.A1(_00706_),
    .A2(_00707_),
    .ZN(_00708_));
 AOI21_X1 _23839_ (.A(_00699_),
    .B1(_21401_),
    .B2(_00708_),
    .ZN(_00709_));
 OAI21_X1 _23840_ (.A(_00678_),
    .B1(_00698_),
    .B2(_00709_),
    .ZN(_00710_));
 NAND3_X1 _23841_ (.A1(_13237_),
    .A2(_00693_),
    .A3(_00620_),
    .ZN(_00711_));
 NOR2_X1 _23842_ (.A1(_13146_),
    .A2(_13241_),
    .ZN(_00712_));
 OAI21_X1 _23843_ (.A(_00636_),
    .B1(_00712_),
    .B2(_00687_),
    .ZN(_00713_));
 OAI21_X1 _23844_ (.A(_00711_),
    .B1(_00713_),
    .B2(_00653_),
    .ZN(_00714_));
 NAND3_X1 _23845_ (.A1(_00699_),
    .A2(_00673_),
    .A3(_00714_),
    .ZN(_00715_));
 OAI21_X1 _23846_ (.A(_13241_),
    .B1(_13229_),
    .B2(_00687_),
    .ZN(_00716_));
 OAI21_X1 _23847_ (.A(_21401_),
    .B1(_00716_),
    .B2(_00653_),
    .ZN(_00717_));
 NAND4_X1 _23848_ (.A1(_00674_),
    .A2(_00654_),
    .A3(_13226_),
    .A4(_13241_),
    .ZN(_00718_));
 NAND2_X1 _23849_ (.A1(_13226_),
    .A2(_00620_),
    .ZN(_00719_));
 NOR2_X1 _23850_ (.A1(_13142_),
    .A2(_13231_),
    .ZN(_00720_));
 OAI221_X2 _23851_ (.A(_00718_),
    .B1(_00719_),
    .B2(_00639_),
    .C1(_13217_),
    .C2(_00720_),
    .ZN(_00721_));
 OAI21_X1 _23852_ (.A(_00717_),
    .B1(_00721_),
    .B2(_21401_),
    .ZN(_00722_));
 OAI21_X1 _23853_ (.A(_00715_),
    .B1(_00722_),
    .B2(_00699_),
    .ZN(_00723_));
 OAI21_X2 _23854_ (.A(_00710_),
    .B1(_00723_),
    .B2(_00678_),
    .ZN(_00724_));
 AOI21_X4 _23855_ (.A(_00684_),
    .B1(_00724_),
    .B2(_00674_),
    .ZN(_00725_));
 NAND2_X2 _23856_ (.A1(_00621_),
    .A2(_00645_),
    .ZN(_00726_));
 NAND2_X1 _23857_ (.A1(_13119_),
    .A2(_13235_),
    .ZN(_00727_));
 NAND2_X1 _23858_ (.A1(_13097_),
    .A2(_00650_),
    .ZN(_00728_));
 MUX2_X2 _23859_ (.A(_00727_),
    .B(_00728_),
    .S(_13140_),
    .Z(_00729_));
 OAI21_X1 _23860_ (.A(_00636_),
    .B1(_13229_),
    .B2(_00729_),
    .ZN(_00730_));
 OAI21_X1 _23861_ (.A(_13229_),
    .B1(_13195_),
    .B2(_00687_),
    .ZN(_00731_));
 OAI21_X1 _23862_ (.A(_00730_),
    .B1(_00731_),
    .B2(_00653_),
    .ZN(_00732_));
 OAI21_X1 _23863_ (.A(_13149_),
    .B1(_13232_),
    .B2(_13142_),
    .ZN(_00733_));
 NOR2_X1 _23864_ (.A1(_13149_),
    .A2(_00693_),
    .ZN(_00734_));
 AOI221_X2 _23865_ (.A(_13221_),
    .B1(_00734_),
    .B2(_00674_),
    .C1(_13142_),
    .C2(_13226_),
    .ZN(_00735_));
 NOR2_X1 _23866_ (.A1(_21401_),
    .A2(_00735_),
    .ZN(_00736_));
 AOI221_X1 _23867_ (.A(_00699_),
    .B1(_21401_),
    .B2(_00732_),
    .C1(_00733_),
    .C2(_00736_),
    .ZN(_00737_));
 NOR2_X1 _23868_ (.A1(_00726_),
    .A2(_00737_),
    .ZN(_00738_));
 NOR3_X1 _23869_ (.A1(_13142_),
    .A2(_13241_),
    .A3(_00673_),
    .ZN(_00739_));
 OAI21_X1 _23870_ (.A(_13156_),
    .B1(_13232_),
    .B2(_13142_),
    .ZN(_00740_));
 OR2_X1 _23871_ (.A1(_13156_),
    .A2(_00693_),
    .ZN(_00741_));
 OAI221_X2 _23872_ (.A(_13217_),
    .B1(_00741_),
    .B2(_00653_),
    .C1(_00729_),
    .C2(_13156_),
    .ZN(_00742_));
 NAND2_X1 _23873_ (.A1(_00740_),
    .A2(_00742_),
    .ZN(_00743_));
 AOI21_X1 _23874_ (.A(_00739_),
    .B1(_00743_),
    .B2(_00673_),
    .ZN(_00744_));
 OAI21_X1 _23875_ (.A(_00738_),
    .B1(_00744_),
    .B2(_00649_),
    .ZN(_00745_));
 MUX2_X1 _23876_ (.A(_00674_),
    .B(_00654_),
    .S(_00624_),
    .Z(_00746_));
 AOI211_X2 _23877_ (.A(_00648_),
    .B(_13115_),
    .C1(_13140_),
    .C2(_13133_),
    .ZN(_00747_));
 AND2_X1 _23878_ (.A1(_13159_),
    .A2(_00747_),
    .ZN(_00748_));
 OAI21_X1 _23879_ (.A(_00748_),
    .B1(_13232_),
    .B2(_13142_),
    .ZN(_00749_));
 AOI211_X2 _23880_ (.A(_00647_),
    .B(_00653_),
    .C1(_00687_),
    .C2(_00626_),
    .ZN(_00750_));
 NAND2_X1 _23881_ (.A1(_00654_),
    .A2(_13230_),
    .ZN(_00751_));
 NAND3_X1 _23882_ (.A1(_13173_),
    .A2(_13184_),
    .A3(_13231_),
    .ZN(_00752_));
 OAI221_X2 _23883_ (.A(_00750_),
    .B1(_00751_),
    .B2(_00630_),
    .C1(_13160_),
    .C2(_00752_),
    .ZN(_00753_));
 NAND4_X1 _23884_ (.A1(_00654_),
    .A2(_13241_),
    .A3(_13223_),
    .A4(_00747_),
    .ZN(_00754_));
 NAND3_X1 _23885_ (.A1(_00729_),
    .A2(_13223_),
    .A3(_00747_),
    .ZN(_00755_));
 NAND3_X2 _23886_ (.A1(_13173_),
    .A2(_13184_),
    .A3(_00638_),
    .ZN(_00756_));
 MUX2_X1 _23887_ (.A(_00754_),
    .B(_00755_),
    .S(_00756_),
    .Z(_00757_));
 AND3_X1 _23888_ (.A1(_00749_),
    .A2(_00753_),
    .A3(_00757_),
    .ZN(_00758_));
 NAND2_X1 _23889_ (.A1(_21401_),
    .A2(_00758_),
    .ZN(_00759_));
 NAND2_X1 _23890_ (.A1(_00672_),
    .A2(_00673_),
    .ZN(_00760_));
 NAND4_X1 _23891_ (.A1(_00683_),
    .A2(_00678_),
    .A3(_00759_),
    .A4(_00760_),
    .ZN(_00761_));
 NAND3_X1 _23892_ (.A1(_00745_),
    .A2(_00746_),
    .A3(_00761_),
    .ZN(_00762_));
 AND4_X1 _23893_ (.A1(_00649_),
    .A2(_00635_),
    .A3(_00645_),
    .A4(_00708_),
    .ZN(_00763_));
 NOR2_X1 _23894_ (.A1(_13254_),
    .A2(_00642_),
    .ZN(_00764_));
 OAI21_X1 _23895_ (.A(_00637_),
    .B1(_00632_),
    .B2(_00764_),
    .ZN(_00765_));
 OAI21_X2 _23896_ (.A(_00675_),
    .B1(_00765_),
    .B2(_00756_),
    .ZN(_00766_));
 NOR3_X1 _23897_ (.A1(_00649_),
    .A2(_00660_),
    .A3(_00766_),
    .ZN(_00767_));
 MUX2_X1 _23898_ (.A(_13226_),
    .B(_13221_),
    .S(_00623_),
    .Z(_00768_));
 AOI221_X2 _23899_ (.A(_00763_),
    .B1(_00767_),
    .B2(_00697_),
    .C1(_00660_),
    .C2(_00768_),
    .ZN(_00769_));
 INV_X1 _23900_ (.A(_00769_),
    .ZN(_00770_));
 OAI21_X1 _23901_ (.A(_00632_),
    .B1(_13159_),
    .B2(_00622_),
    .ZN(_00771_));
 AND2_X1 _23902_ (.A1(_21401_),
    .A2(_00771_),
    .ZN(_00772_));
 NAND4_X2 _23903_ (.A1(_00749_),
    .A2(_00753_),
    .A3(_00757_),
    .A4(_00772_),
    .ZN(_00773_));
 OAI21_X1 _23904_ (.A(_00771_),
    .B1(_00766_),
    .B2(_00632_),
    .ZN(_00774_));
 NAND3_X1 _23905_ (.A1(_00672_),
    .A2(_00616_),
    .A3(_00771_),
    .ZN(_00775_));
 NAND3_X2 _23906_ (.A1(_00622_),
    .A2(_00689_),
    .A3(_00660_),
    .ZN(_00776_));
 NAND4_X4 _23907_ (.A1(_00773_),
    .A2(_00774_),
    .A3(_00775_),
    .A4(_00776_),
    .ZN(_00777_));
 NOR3_X2 _23908_ (.A1(_00624_),
    .A2(_13159_),
    .A3(_00621_),
    .ZN(_00778_));
 OAI21_X1 _23909_ (.A(_00660_),
    .B1(_13223_),
    .B2(_00658_),
    .ZN(_00779_));
 AND2_X1 _23910_ (.A1(_00635_),
    .A2(_00645_),
    .ZN(_00780_));
 MUX2_X1 _23911_ (.A(_00685_),
    .B(_00708_),
    .S(_00699_),
    .Z(_00781_));
 NAND2_X1 _23912_ (.A1(_00780_),
    .A2(_00781_),
    .ZN(_00782_));
 AOI211_X2 _23913_ (.A(_00777_),
    .B(_00778_),
    .C1(_00779_),
    .C2(_00782_),
    .ZN(_00783_));
 AND3_X1 _23914_ (.A1(_21383_),
    .A2(_00770_),
    .A3(_00783_),
    .ZN(_00784_));
 NOR2_X1 _23915_ (.A1(_00624_),
    .A2(_00687_),
    .ZN(_00785_));
 NOR2_X1 _23916_ (.A1(_00658_),
    .A2(_13241_),
    .ZN(_00786_));
 NOR3_X1 _23917_ (.A1(_00686_),
    .A2(_00688_),
    .A3(_00695_),
    .ZN(_00787_));
 NAND2_X1 _23918_ (.A1(_00673_),
    .A2(_00787_),
    .ZN(_00788_));
 OAI21_X1 _23919_ (.A(_00788_),
    .B1(_00714_),
    .B2(_00673_),
    .ZN(_00789_));
 OAI33_X1 _23920_ (.A1(_00621_),
    .A2(_00785_),
    .A3(_00786_),
    .B1(_00789_),
    .B2(_00726_),
    .B3(_00699_),
    .ZN(_00790_));
 NOR3_X1 _23921_ (.A1(_00649_),
    .A2(_00726_),
    .A3(_00722_),
    .ZN(_00791_));
 AND3_X1 _23922_ (.A1(_00635_),
    .A2(_00678_),
    .A3(_00781_),
    .ZN(_00792_));
 OR3_X2 _23923_ (.A1(_00790_),
    .A2(_00791_),
    .A3(_00792_),
    .ZN(_00793_));
 NOR2_X1 _23924_ (.A1(_00622_),
    .A2(_13156_),
    .ZN(_00794_));
 NOR2_X1 _23925_ (.A1(_00623_),
    .A2(_13260_),
    .ZN(_00795_));
 OAI21_X1 _23926_ (.A(_00620_),
    .B1(_00616_),
    .B2(_00672_),
    .ZN(_00796_));
 OAI33_X1 _23927_ (.A1(_00621_),
    .A2(_00794_),
    .A3(_00795_),
    .B1(_00796_),
    .B2(_00677_),
    .B3(_13142_),
    .ZN(_00797_));
 NOR3_X2 _23928_ (.A1(_00660_),
    .A2(_21401_),
    .A3(_00766_),
    .ZN(_00798_));
 NOR3_X1 _23929_ (.A1(_00699_),
    .A2(_00653_),
    .A3(_00735_),
    .ZN(_00799_));
 AND2_X1 _23930_ (.A1(_00747_),
    .A2(_00742_),
    .ZN(_00800_));
 AOI22_X2 _23931_ (.A1(_00733_),
    .A2(_00799_),
    .B1(_00800_),
    .B2(_00740_),
    .ZN(_00801_));
 AOI221_X2 _23932_ (.A(_00797_),
    .B1(_00798_),
    .B2(_00758_),
    .C1(_00801_),
    .C2(_00780_),
    .ZN(_00802_));
 MUX2_X1 _23933_ (.A(_13149_),
    .B(_13217_),
    .S(_00658_),
    .Z(_00803_));
 AND2_X1 _23934_ (.A1(_00647_),
    .A2(_00735_),
    .ZN(_00804_));
 NOR3_X1 _23935_ (.A1(_00648_),
    .A2(_13226_),
    .A3(_00752_),
    .ZN(_00805_));
 NOR2_X1 _23936_ (.A1(_00647_),
    .A2(_13159_),
    .ZN(_00806_));
 AND2_X1 _23937_ (.A1(_13232_),
    .A2(_00806_),
    .ZN(_00807_));
 NAND3_X1 _23938_ (.A1(_00648_),
    .A2(_00729_),
    .A3(_00659_),
    .ZN(_00808_));
 AOI21_X1 _23939_ (.A(_00806_),
    .B1(_13149_),
    .B2(_00647_),
    .ZN(_00809_));
 OAI22_X1 _23940_ (.A1(_13232_),
    .A2(_00808_),
    .B1(_00809_),
    .B2(_00729_),
    .ZN(_00810_));
 OR4_X2 _23941_ (.A1(_00804_),
    .A2(_00805_),
    .A3(_00807_),
    .A4(_00810_),
    .ZN(_00811_));
 NAND3_X2 _23942_ (.A1(_00621_),
    .A2(_00616_),
    .A3(_00645_),
    .ZN(_00812_));
 OAI222_X2 _23943_ (.A1(_00621_),
    .A2(_00803_),
    .B1(_00811_),
    .B2(_00646_),
    .C1(_00666_),
    .C2(_00812_),
    .ZN(_00813_));
 NAND3_X1 _23944_ (.A1(_00673_),
    .A2(_00706_),
    .A3(_00707_),
    .ZN(_00814_));
 OAI211_X2 _23945_ (.A(_00699_),
    .B(_00814_),
    .C1(_00721_),
    .C2(_00673_),
    .ZN(_00815_));
 OAI21_X1 _23946_ (.A(_00616_),
    .B1(_00655_),
    .B2(_00653_),
    .ZN(_00816_));
 OAI211_X2 _23947_ (.A(_00649_),
    .B(_00816_),
    .C1(_00696_),
    .C2(_00673_),
    .ZN(_00817_));
 AOI21_X2 _23948_ (.A(_00726_),
    .B1(_00815_),
    .B2(_00817_),
    .ZN(_00818_));
 MUX2_X1 _23949_ (.A(_13156_),
    .B(_13217_),
    .S(_00624_),
    .Z(_00819_));
 NOR2_X1 _23950_ (.A1(_00621_),
    .A2(_00819_),
    .ZN(_00820_));
 OAI211_X2 _23951_ (.A(_00802_),
    .B(_00813_),
    .C1(_00818_),
    .C2(_00820_),
    .ZN(_00821_));
 NOR2_X1 _23952_ (.A1(_00658_),
    .A2(_13229_),
    .ZN(_00822_));
 NOR2_X1 _23953_ (.A1(_00624_),
    .A2(_13241_),
    .ZN(_00823_));
 NOR2_X1 _23954_ (.A1(_13239_),
    .A2(_00643_),
    .ZN(_00824_));
 OAI21_X1 _23955_ (.A(_00824_),
    .B1(_13232_),
    .B2(_13142_),
    .ZN(_00825_));
 MUX2_X1 _23956_ (.A(_13250_),
    .B(_00825_),
    .S(_13233_),
    .Z(_00826_));
 NAND2_X1 _23957_ (.A1(_00637_),
    .A2(_00620_),
    .ZN(_00827_));
 OAI33_X1 _23958_ (.A1(_00621_),
    .A2(_00822_),
    .A3(_00823_),
    .B1(_00826_),
    .B2(_00827_),
    .B3(_00666_),
    .ZN(_00828_));
 NOR2_X1 _23959_ (.A1(_00812_),
    .A2(_00811_),
    .ZN(_00829_));
 INV_X1 _23960_ (.A(_00732_),
    .ZN(_00830_));
 AOI21_X1 _23961_ (.A(_00646_),
    .B1(_00830_),
    .B2(_00699_),
    .ZN(_00831_));
 NAND2_X1 _23962_ (.A1(_00649_),
    .A2(_00743_),
    .ZN(_00832_));
 AOI211_X2 _23963_ (.A(_00828_),
    .B(_00829_),
    .C1(_00831_),
    .C2(_00832_),
    .ZN(_00833_));
 OAI21_X1 _23964_ (.A(_00635_),
    .B1(_00721_),
    .B2(_00699_),
    .ZN(_00834_));
 OR3_X1 _23965_ (.A1(_00632_),
    .A2(_00677_),
    .A3(_00655_),
    .ZN(_00835_));
 NOR2_X1 _23966_ (.A1(_00649_),
    .A2(_00714_),
    .ZN(_00836_));
 AOI21_X1 _23967_ (.A(_00834_),
    .B1(_00835_),
    .B2(_00836_),
    .ZN(_00837_));
 MUX2_X1 _23968_ (.A(_00696_),
    .B(_00708_),
    .S(_00649_),
    .Z(_00838_));
 MUX2_X1 _23969_ (.A(_13229_),
    .B(_00636_),
    .S(_00624_),
    .Z(_00839_));
 AOI221_X2 _23970_ (.A(_00837_),
    .B1(_00838_),
    .B2(_00798_),
    .C1(_00660_),
    .C2(_00839_),
    .ZN(_00840_));
 NOR3_X1 _23971_ (.A1(_00821_),
    .A2(_00833_),
    .A3(_00840_),
    .ZN(_00841_));
 NAND4_X2 _23972_ (.A1(_00762_),
    .A2(_00784_),
    .A3(_00793_),
    .A4(_00841_),
    .ZN(_00842_));
 XOR2_X2 _23973_ (.A(_00725_),
    .B(_00842_),
    .Z(_00843_));
 MUX2_X1 _23974_ (.A(_00671_),
    .B(_00682_),
    .S(_00843_),
    .Z(_00844_));
 OR2_X2 _23975_ (.A1(_00668_),
    .A2(_12835_),
    .ZN(_00845_));
 OAI21_X1 _23976_ (.A(_00670_),
    .B1(_00844_),
    .B2(_00845_),
    .ZN(_00048_));
 AOI22_X1 _23977_ (.A1(\g_reduce0[14].adder.b[1] ),
    .A2(_00668_),
    .B1(_00669_),
    .B2(\g_reduce0[14].adder.a[1] ),
    .ZN(_00846_));
 INV_X1 _23978_ (.A(_21385_),
    .ZN(_00847_));
 XNOR2_X1 _23979_ (.A(_00847_),
    .B(_00777_),
    .ZN(_00848_));
 MUX2_X1 _23980_ (.A(_00848_),
    .B(_00671_),
    .S(_00843_),
    .Z(_00849_));
 OAI21_X1 _23981_ (.A(_00846_),
    .B1(_00849_),
    .B2(_00845_),
    .ZN(_00055_));
 AOI21_X1 _23982_ (.A(_00770_),
    .B1(_00783_),
    .B2(_21383_),
    .ZN(_00850_));
 NOR2_X1 _23983_ (.A1(_00784_),
    .A2(_00850_),
    .ZN(_00851_));
 NOR3_X1 _23984_ (.A1(_00845_),
    .A2(_00843_),
    .A3(_00851_),
    .ZN(_00852_));
 NOR2_X2 _23985_ (.A1(_00668_),
    .A2(_12835_),
    .ZN(_00853_));
 AND3_X1 _23986_ (.A1(_00853_),
    .A2(_00843_),
    .A3(_00848_),
    .ZN(_00854_));
 NAND2_X1 _23987_ (.A1(_12832_),
    .A2(_12836_),
    .ZN(_00855_));
 OAI22_X1 _23988_ (.A1(\g_reduce0[14].adder.b[2] ),
    .A2(_12833_),
    .B1(_00855_),
    .B2(\g_reduce0[14].adder.a[2] ),
    .ZN(_00856_));
 NOR3_X1 _23989_ (.A1(_00852_),
    .A2(_00854_),
    .A3(_00856_),
    .ZN(_00056_));
 NOR2_X1 _23990_ (.A1(_00845_),
    .A2(_00851_),
    .ZN(_00857_));
 NAND2_X1 _23991_ (.A1(_00843_),
    .A2(_00857_),
    .ZN(_00858_));
 NOR3_X2 _23992_ (.A1(_00847_),
    .A2(_00777_),
    .A3(_00769_),
    .ZN(_00859_));
 XNOR2_X1 _23993_ (.A(_00813_),
    .B(_00859_),
    .ZN(_00860_));
 NAND2_X1 _23994_ (.A1(_00853_),
    .A2(_00860_),
    .ZN(_00861_));
 OAI21_X1 _23995_ (.A(_00858_),
    .B1(_00861_),
    .B2(_00843_),
    .ZN(_00862_));
 OAI22_X1 _23996_ (.A1(\g_reduce0[14].adder.b[3] ),
    .A2(_12833_),
    .B1(_00855_),
    .B2(\g_reduce0[14].adder.a[3] ),
    .ZN(_00863_));
 NOR2_X1 _23997_ (.A1(_00862_),
    .A2(_00863_),
    .ZN(_00057_));
 AOI22_X1 _23998_ (.A1(\g_reduce0[14].adder.b[4] ),
    .A2(_00668_),
    .B1(_00669_),
    .B2(\g_reduce0[14].adder.a[4] ),
    .ZN(_00864_));
 NOR2_X1 _23999_ (.A1(_00820_),
    .A2(_00818_),
    .ZN(_00865_));
 NAND3_X2 _24000_ (.A1(_21383_),
    .A2(_00770_),
    .A3(_00783_),
    .ZN(_00866_));
 NOR2_X1 _24001_ (.A1(_00646_),
    .A2(_00811_),
    .ZN(_00867_));
 OAI22_X1 _24002_ (.A1(_00666_),
    .A2(_00812_),
    .B1(_00803_),
    .B2(_00683_),
    .ZN(_00868_));
 NOR2_X1 _24003_ (.A1(_00867_),
    .A2(_00868_),
    .ZN(_00869_));
 NOR2_X1 _24004_ (.A1(_00866_),
    .A2(_00869_),
    .ZN(_00870_));
 XOR2_X1 _24005_ (.A(_00865_),
    .B(_00870_),
    .Z(_00871_));
 MUX2_X1 _24006_ (.A(_00871_),
    .B(_00860_),
    .S(_00843_),
    .Z(_00872_));
 OAI21_X1 _24007_ (.A(_00864_),
    .B1(_00872_),
    .B2(_00845_),
    .ZN(_00058_));
 OAI22_X1 _24008_ (.A1(\g_reduce0[14].adder.b[5] ),
    .A2(_12833_),
    .B1(_00855_),
    .B2(\g_reduce0[14].adder.a[5] ),
    .ZN(_00873_));
 OR3_X1 _24009_ (.A1(_00847_),
    .A2(_00777_),
    .A3(_00769_),
    .ZN(_00874_));
 NOR3_X1 _24010_ (.A1(_00865_),
    .A2(_00869_),
    .A3(_00874_),
    .ZN(_00875_));
 XNOR2_X1 _24011_ (.A(_00802_),
    .B(_00875_),
    .ZN(_00876_));
 MUX2_X1 _24012_ (.A(_00876_),
    .B(_00871_),
    .S(_00843_),
    .Z(_00877_));
 AOI21_X1 _24013_ (.A(_00873_),
    .B1(_00877_),
    .B2(_00853_),
    .ZN(_00059_));
 OAI22_X1 _24014_ (.A1(\g_reduce0[14].adder.b[6] ),
    .A2(_12833_),
    .B1(_00855_),
    .B2(\g_reduce0[14].adder.a[6] ),
    .ZN(_00878_));
 INV_X1 _24015_ (.A(_00762_),
    .ZN(_00879_));
 NAND2_X1 _24016_ (.A1(_00793_),
    .A2(_00841_),
    .ZN(_00880_));
 NOR3_X1 _24017_ (.A1(_00879_),
    .A2(_00866_),
    .A3(_00880_),
    .ZN(_00881_));
 OR2_X1 _24018_ (.A1(_00881_),
    .A2(_00876_),
    .ZN(_00882_));
 NOR2_X1 _24019_ (.A1(_00866_),
    .A2(_00821_),
    .ZN(_00883_));
 XNOR2_X1 _24020_ (.A(_00840_),
    .B(_00883_),
    .ZN(_00884_));
 NOR2_X1 _24021_ (.A1(_00842_),
    .A2(_00859_),
    .ZN(_00885_));
 NOR2_X1 _24022_ (.A1(_00884_),
    .A2(_00885_),
    .ZN(_00886_));
 MUX2_X1 _24023_ (.A(_00882_),
    .B(_00886_),
    .S(_00725_),
    .Z(_00887_));
 AOI21_X1 _24024_ (.A(_00878_),
    .B1(_00887_),
    .B2(_00853_),
    .ZN(_00060_));
 AOI22_X1 _24025_ (.A1(\g_reduce0[14].adder.b[7] ),
    .A2(_00668_),
    .B1(_00669_),
    .B2(\g_reduce0[14].adder.a[7] ),
    .ZN(_00888_));
 OR2_X1 _24026_ (.A1(_00821_),
    .A2(_00840_),
    .ZN(_00889_));
 OR3_X1 _24027_ (.A1(_00833_),
    .A2(_00889_),
    .A3(_00874_),
    .ZN(_00890_));
 OAI21_X1 _24028_ (.A(_00833_),
    .B1(_00889_),
    .B2(_00874_),
    .ZN(_00891_));
 NAND3_X1 _24029_ (.A1(_00842_),
    .A2(_00890_),
    .A3(_00891_),
    .ZN(_00892_));
 MUX2_X1 _24030_ (.A(_00886_),
    .B(_00892_),
    .S(_00725_),
    .Z(_00893_));
 OAI21_X1 _24031_ (.A(_00888_),
    .B1(_00893_),
    .B2(_00845_),
    .ZN(_00061_));
 NAND2_X1 _24032_ (.A1(_00853_),
    .A2(_00725_),
    .ZN(_00894_));
 NAND2_X1 _24033_ (.A1(_00784_),
    .A2(_00841_),
    .ZN(_00895_));
 XNOR2_X1 _24034_ (.A(_00793_),
    .B(_00895_),
    .ZN(_00896_));
 NOR3_X1 _24035_ (.A1(_00885_),
    .A2(_00894_),
    .A3(_00896_),
    .ZN(_00897_));
 NOR2_X1 _24036_ (.A1(_12835_),
    .A2(_00725_),
    .ZN(_00898_));
 INV_X1 _24037_ (.A(\g_reduce0[14].adder.a[8] ),
    .ZN(_00899_));
 AOI221_X2 _24038_ (.A(_00668_),
    .B1(_00892_),
    .B2(_00898_),
    .C1(_12836_),
    .C2(_00899_),
    .ZN(_00900_));
 AOI21_X1 _24039_ (.A(_00900_),
    .B1(_00668_),
    .B2(\g_reduce0[14].adder.b[8] ),
    .ZN(_00901_));
 NOR2_X1 _24040_ (.A1(_00897_),
    .A2(_00901_),
    .ZN(_00062_));
 AOI22_X1 _24041_ (.A1(\g_reduce0[14].adder.b[9] ),
    .A2(_00668_),
    .B1(_00669_),
    .B2(\g_reduce0[14].adder.a[9] ),
    .ZN(_00902_));
 AOI21_X1 _24042_ (.A(_00880_),
    .B1(_00874_),
    .B2(_00866_),
    .ZN(_00903_));
 NAND2_X1 _24043_ (.A1(_00879_),
    .A2(_00859_),
    .ZN(_00904_));
 OAI221_X1 _24044_ (.A(_00725_),
    .B1(_00879_),
    .B2(_00903_),
    .C1(_00904_),
    .C2(_00880_),
    .ZN(_00905_));
 NAND2_X1 _24045_ (.A1(_00853_),
    .A2(_00905_),
    .ZN(_00906_));
 NOR3_X1 _24046_ (.A1(_00725_),
    .A2(_00885_),
    .A3(_00896_),
    .ZN(_00907_));
 OAI21_X1 _24047_ (.A(_00902_),
    .B1(_00906_),
    .B2(_00907_),
    .ZN(_00063_));
 INV_X1 _24048_ (.A(_21387_),
    .ZN(_21393_));
 MUX2_X1 _24049_ (.A(_21392_),
    .B(\g_reduce0[14].adder.a[10] ),
    .S(_12836_),
    .Z(_00908_));
 MUX2_X1 _24050_ (.A(\g_reduce0[14].adder.b[10] ),
    .B(_00908_),
    .S(_12833_),
    .Z(_00049_));
 MUX2_X1 _24051_ (.A(_21400_),
    .B(_12829_),
    .S(_12836_),
    .Z(_00909_));
 MUX2_X1 _24052_ (.A(\g_reduce0[14].adder.b[11] ),
    .B(_00909_),
    .S(_12833_),
    .Z(_00050_));
 MUX2_X1 _24053_ (.A(_21265_),
    .B(_00500_),
    .S(_12877_),
    .Z(_00910_));
 NAND2_X1 _24054_ (.A1(_00658_),
    .A2(_21394_),
    .ZN(_00911_));
 XOR2_X1 _24055_ (.A(_00910_),
    .B(_00911_),
    .Z(_00912_));
 XOR2_X1 _24056_ (.A(_14085_),
    .B(_21404_),
    .Z(_00913_));
 MUX2_X1 _24057_ (.A(_00912_),
    .B(_00913_),
    .S(_00683_),
    .Z(_00914_));
 XOR2_X1 _24058_ (.A(_21399_),
    .B(_00914_),
    .Z(_00915_));
 MUX2_X1 _24059_ (.A(_00915_),
    .B(\g_reduce0[14].adder.a[12] ),
    .S(_12836_),
    .Z(_00916_));
 MUX2_X1 _24060_ (.A(\g_reduce0[14].adder.b[12] ),
    .B(_00916_),
    .S(_12833_),
    .Z(_00051_));
 INV_X1 _24061_ (.A(_14087_),
    .ZN(_14084_));
 MUX2_X1 _24062_ (.A(_21262_),
    .B(_00503_),
    .S(_12877_),
    .Z(_00917_));
 MUX2_X1 _24063_ (.A(_21268_),
    .B(_00495_),
    .S(_12877_),
    .Z(_00918_));
 NOR4_X1 _24064_ (.A1(_00624_),
    .A2(_21387_),
    .A3(_00910_),
    .A4(_00918_),
    .ZN(_00919_));
 XNOR2_X1 _24065_ (.A(_00917_),
    .B(_00919_),
    .ZN(_00920_));
 INV_X1 _24066_ (.A(_21396_),
    .ZN(_00921_));
 INV_X1 _24067_ (.A(_21397_),
    .ZN(_00922_));
 OAI21_X1 _24068_ (.A(_00921_),
    .B1(_00922_),
    .B2(_14087_),
    .ZN(_00923_));
 AOI21_X1 _24069_ (.A(_21403_),
    .B1(_00923_),
    .B2(_21404_),
    .ZN(_00924_));
 XNOR2_X1 _24070_ (.A(_21408_),
    .B(_00924_),
    .ZN(_00925_));
 MUX2_X1 _24071_ (.A(_00920_),
    .B(_00925_),
    .S(_00683_),
    .Z(_00926_));
 NAND2_X1 _24072_ (.A1(_00658_),
    .A2(_21395_),
    .ZN(_00927_));
 OAI21_X1 _24073_ (.A(_00927_),
    .B1(_00918_),
    .B2(_00658_),
    .ZN(_00928_));
 MUX2_X1 _24074_ (.A(_14086_),
    .B(_00928_),
    .S(_00660_),
    .Z(_21398_));
 NAND3_X1 _24075_ (.A1(_21391_),
    .A2(_00914_),
    .A3(_21398_),
    .ZN(_00929_));
 XNOR2_X1 _24076_ (.A(_00926_),
    .B(_00929_),
    .ZN(_00930_));
 MUX2_X1 _24077_ (.A(_00930_),
    .B(\g_reduce0[14].adder.a[13] ),
    .S(_12836_),
    .Z(_00931_));
 MUX2_X1 _24078_ (.A(\g_reduce0[14].adder.b[13] ),
    .B(_00931_),
    .S(_12833_),
    .Z(_00052_));
 AND2_X1 _24079_ (.A1(\g_reduce0[14].adder.b[14] ),
    .A2(_12849_),
    .ZN(_00932_));
 NOR4_X1 _24080_ (.A1(_00683_),
    .A2(_00910_),
    .A3(_00911_),
    .A4(_00917_),
    .ZN(_00933_));
 AOI21_X1 _24081_ (.A(_21403_),
    .B1(_21404_),
    .B2(_14085_),
    .ZN(_00934_));
 INV_X1 _24082_ (.A(_00934_),
    .ZN(_00935_));
 AOI21_X1 _24083_ (.A(_21407_),
    .B1(_00935_),
    .B2(_21408_),
    .ZN(_00936_));
 AOI21_X1 _24084_ (.A(_00933_),
    .B1(_00936_),
    .B2(_00683_),
    .ZN(_00937_));
 NAND3_X1 _24085_ (.A1(_21399_),
    .A2(_00914_),
    .A3(_00926_),
    .ZN(_00938_));
 XOR2_X2 _24086_ (.A(_00937_),
    .B(_00938_),
    .Z(_00939_));
 MUX2_X1 _24087_ (.A(_12881_),
    .B(_00932_),
    .S(_00939_),
    .Z(_00940_));
 NOR2_X1 _24088_ (.A1(_12836_),
    .A2(_00940_),
    .ZN(_00941_));
 NOR3_X1 _24089_ (.A1(_12830_),
    .A2(_00668_),
    .A3(_00941_),
    .ZN(_00942_));
 OR2_X1 _24090_ (.A1(\g_reduce0[14].adder.b[14] ),
    .A2(_12881_),
    .ZN(_00943_));
 NAND2_X1 _24091_ (.A1(_12830_),
    .A2(_00943_),
    .ZN(_00944_));
 MUX2_X1 _24092_ (.A(_00943_),
    .B(_00944_),
    .S(_00939_),
    .Z(_00945_));
 OAI22_X1 _24093_ (.A1(\g_reduce0[14].adder.b[14] ),
    .A2(_12833_),
    .B1(_12836_),
    .B2(_00945_),
    .ZN(_00946_));
 NOR2_X1 _24094_ (.A1(_00942_),
    .A2(_00946_),
    .ZN(_00053_));
 CLKBUF_X2 _24095_ (.A(\g_reduce0[2].adder.b[15] ),
    .Z(_00947_));
 CLKBUF_X2 _24096_ (.A(\g_reduce0[2].adder.a[15] ),
    .Z(_00948_));
 OR3_X1 _24097_ (.A1(\g_reduce0[2].adder.a[11] ),
    .A2(\g_reduce0[2].adder.a[10] ),
    .A3(\g_reduce0[2].adder.a[13] ),
    .ZN(_00949_));
 NOR3_X2 _24098_ (.A1(\g_reduce0[2].adder.a[12] ),
    .A2(\g_reduce0[2].adder.a[14] ),
    .A3(_00949_),
    .ZN(_00950_));
 CLKBUF_X3 _24099_ (.A(_00950_),
    .Z(_00951_));
 BUF_X2 _24100_ (.A(\g_reduce0[2].adder.b[11] ),
    .Z(_00952_));
 BUF_X2 _24101_ (.A(\g_reduce0[2].adder.b[14] ),
    .Z(_00953_));
 OR2_X1 _24102_ (.A1(\g_reduce0[2].adder.b[10] ),
    .A2(\g_reduce0[2].adder.b[13] ),
    .ZN(_00954_));
 OR4_X1 _24103_ (.A1(_00952_),
    .A2(\g_reduce0[2].adder.b[12] ),
    .A3(_00953_),
    .A4(_00954_),
    .ZN(_00955_));
 BUF_X2 _24104_ (.A(_00955_),
    .Z(_00956_));
 CLKBUF_X3 _24105_ (.A(_00956_),
    .Z(_00957_));
 BUF_X2 _24106_ (.A(_21456_),
    .Z(_00958_));
 INV_X2 _24107_ (.A(_00958_),
    .ZN(_00959_));
 BUF_X2 _24108_ (.A(_21450_),
    .Z(_00960_));
 INV_X4 _24109_ (.A(_00960_),
    .ZN(_00961_));
 INV_X2 _24110_ (.A(_21417_),
    .ZN(_00962_));
 BUF_X2 _24111_ (.A(_21411_),
    .Z(_00963_));
 BUF_X4 _24112_ (.A(_21414_),
    .Z(_00964_));
 NAND2_X4 _24113_ (.A1(_00963_),
    .A2(_00964_),
    .ZN(_00965_));
 NOR4_X1 _24114_ (.A1(_00959_),
    .A2(_00961_),
    .A3(_00962_),
    .A4(_00965_),
    .ZN(_00966_));
 INV_X1 _24115_ (.A(_21455_),
    .ZN(_00967_));
 AOI21_X2 _24116_ (.A(_21410_),
    .B1(_21413_),
    .B2(_00963_),
    .ZN(_00968_));
 OAI21_X2 _24117_ (.A(_00967_),
    .B1(_00968_),
    .B2(_00959_),
    .ZN(_00969_));
 INV_X1 _24118_ (.A(_21416_),
    .ZN(_00970_));
 OAI21_X2 _24119_ (.A(_00970_),
    .B1(_21449_),
    .B2(_00962_),
    .ZN(_00971_));
 NOR2_X2 _24120_ (.A1(_00959_),
    .A2(_00965_),
    .ZN(_00972_));
 AOI21_X4 _24121_ (.A(_00969_),
    .B1(_00971_),
    .B2(_00972_),
    .ZN(_00973_));
 NOR2_X4 _24122_ (.A1(_00966_),
    .A2(_00973_),
    .ZN(_00974_));
 AND4_X2 _24123_ (.A1(_21420_),
    .A2(_21423_),
    .A3(_21426_),
    .A4(_21429_),
    .ZN(_00975_));
 AND4_X1 _24124_ (.A1(_21432_),
    .A2(_21435_),
    .A3(_21438_),
    .A4(_21441_),
    .ZN(_00976_));
 NAND4_X4 _24125_ (.A1(_21444_),
    .A2(_21447_),
    .A3(_00975_),
    .A4(_00976_),
    .ZN(_00977_));
 INV_X1 _24126_ (.A(_00977_),
    .ZN(_00978_));
 AOI21_X1 _24127_ (.A(_21431_),
    .B1(_21434_),
    .B2(_21432_),
    .ZN(_00979_));
 NAND2_X1 _24128_ (.A1(_21432_),
    .A2(_21435_),
    .ZN(_00980_));
 AOI21_X1 _24129_ (.A(_21437_),
    .B1(_21438_),
    .B2(_21440_),
    .ZN(_00981_));
 OAI21_X2 _24130_ (.A(_00979_),
    .B1(_00980_),
    .B2(_00981_),
    .ZN(_00982_));
 NAND2_X4 _24131_ (.A1(_00975_),
    .A2(_00982_),
    .ZN(_00983_));
 INV_X1 _24132_ (.A(_21443_),
    .ZN(_00984_));
 INV_X1 _24133_ (.A(_21444_),
    .ZN(_00985_));
 OAI21_X1 _24134_ (.A(_00984_),
    .B1(_21446_),
    .B2(_00985_),
    .ZN(_00986_));
 AND2_X1 _24135_ (.A1(_00975_),
    .A2(_00976_),
    .ZN(_00987_));
 INV_X1 _24136_ (.A(_21422_),
    .ZN(_00988_));
 AOI21_X1 _24137_ (.A(_21425_),
    .B1(_21426_),
    .B2(_21428_),
    .ZN(_00989_));
 INV_X1 _24138_ (.A(_21423_),
    .ZN(_00990_));
 OAI21_X1 _24139_ (.A(_00988_),
    .B1(_00989_),
    .B2(_00990_),
    .ZN(_00991_));
 AOI221_X4 _24140_ (.A(_21419_),
    .B1(_00986_),
    .B2(_00987_),
    .C1(_00991_),
    .C2(_21420_),
    .ZN(_00992_));
 AOI21_X4 _24141_ (.A(_00978_),
    .B1(_00983_),
    .B2(_00992_),
    .ZN(_00993_));
 BUF_X1 _24142_ (.A(_00966_),
    .Z(_00994_));
 AOI21_X4 _24143_ (.A(_00974_),
    .B1(_00993_),
    .B2(_00994_),
    .ZN(_00995_));
 AOI21_X2 _24144_ (.A(_00951_),
    .B1(_00957_),
    .B2(_00995_),
    .ZN(_00996_));
 MUX2_X2 _24145_ (.A(_00947_),
    .B(_00948_),
    .S(_00996_),
    .Z(_00070_));
 BUF_X2 _24146_ (.A(_00506_),
    .Z(_00997_));
 NAND3_X2 _24147_ (.A1(_00960_),
    .A2(_21417_),
    .A3(_00972_),
    .ZN(_00998_));
 AND2_X1 _24148_ (.A1(_00963_),
    .A2(_00964_),
    .ZN(_00999_));
 NAND2_X1 _24149_ (.A1(_00958_),
    .A2(_00999_),
    .ZN(_01000_));
 INV_X1 _24150_ (.A(_21449_),
    .ZN(_01001_));
 AOI21_X1 _24151_ (.A(_21416_),
    .B1(_01001_),
    .B2(_21417_),
    .ZN(_01002_));
 OAI221_X1 _24152_ (.A(_00967_),
    .B1(_01000_),
    .B2(_01002_),
    .C1(_00968_),
    .C2(_00959_),
    .ZN(_01003_));
 CLKBUF_X3 _24153_ (.A(_01003_),
    .Z(_01004_));
 NAND2_X2 _24154_ (.A1(_00998_),
    .A2(_01004_),
    .ZN(_01005_));
 INV_X1 _24155_ (.A(_21447_),
    .ZN(_01006_));
 NAND2_X1 _24156_ (.A1(_00975_),
    .A2(_00976_),
    .ZN(_01007_));
 INV_X1 _24157_ (.A(_21419_),
    .ZN(_01008_));
 INV_X1 _24158_ (.A(_21446_),
    .ZN(_01009_));
 AOI21_X1 _24159_ (.A(_21443_),
    .B1(_01009_),
    .B2(_21444_),
    .ZN(_01010_));
 OAI21_X1 _24160_ (.A(_01008_),
    .B1(_01010_),
    .B2(_01007_),
    .ZN(_01011_));
 AND2_X1 _24161_ (.A1(_00975_),
    .A2(_00982_),
    .ZN(_01012_));
 AND2_X1 _24162_ (.A1(_21420_),
    .A2(_00991_),
    .ZN(_01013_));
 OAI33_X1 _24163_ (.A1(_00985_),
    .A2(_01006_),
    .A3(_01007_),
    .B1(_01011_),
    .B2(_01012_),
    .B3(_01013_),
    .ZN(_01014_));
 BUF_X4 _24164_ (.A(_01014_),
    .Z(_01015_));
 BUF_X4 _24165_ (.A(_00998_),
    .Z(_01016_));
 OAI21_X2 _24166_ (.A(_01005_),
    .B1(_01015_),
    .B2(_01016_),
    .ZN(_01017_));
 BUF_X4 _24167_ (.A(_01017_),
    .Z(_01018_));
 MUX2_X2 _24168_ (.A(_00997_),
    .B(_21448_),
    .S(_01018_),
    .Z(_21534_));
 NOR2_X4 _24169_ (.A1(\g_reduce0[2].adder.a[11] ),
    .A2(_21415_),
    .ZN(_01019_));
 OAI211_X4 _24170_ (.A(_01005_),
    .B(_01019_),
    .C1(_01015_),
    .C2(_01016_),
    .ZN(_01020_));
 NOR2_X1 _24171_ (.A1(_00952_),
    .A2(_00509_),
    .ZN(_01021_));
 NAND3_X1 _24172_ (.A1(_00966_),
    .A2(_00977_),
    .A3(_01021_),
    .ZN(_01022_));
 AOI21_X2 _24173_ (.A(_01022_),
    .B1(_00983_),
    .B2(_00992_),
    .ZN(_01023_));
 AND3_X1 _24174_ (.A1(_00998_),
    .A2(_01004_),
    .A3(_01021_),
    .ZN(_01024_));
 NOR3_X4 _24175_ (.A1(_21452_),
    .A2(_01023_),
    .A3(_01024_),
    .ZN(_01025_));
 AOI21_X4 _24176_ (.A(_01000_),
    .B1(_01020_),
    .B2(_01025_),
    .ZN(_01026_));
 NOR2_X1 _24177_ (.A1(\g_reduce0[2].adder.b[13] ),
    .A2(_00517_),
    .ZN(_01027_));
 NAND3_X1 _24178_ (.A1(_00966_),
    .A2(_00977_),
    .A3(_01027_),
    .ZN(_01028_));
 AOI21_X1 _24179_ (.A(_01028_),
    .B1(_00983_),
    .B2(_00992_),
    .ZN(_01029_));
 NOR2_X1 _24180_ (.A1(\g_reduce0[2].adder.a[13] ),
    .A2(_21409_),
    .ZN(_01030_));
 AND2_X1 _24181_ (.A1(_00994_),
    .A2(_01030_),
    .ZN(_01031_));
 MUX2_X1 _24182_ (.A(_01030_),
    .B(_01027_),
    .S(_01004_),
    .Z(_01032_));
 AOI221_X2 _24183_ (.A(_01029_),
    .B1(_01031_),
    .B2(_01015_),
    .C1(_01032_),
    .C2(_01016_),
    .ZN(_01033_));
 NOR2_X2 _24184_ (.A1(_00959_),
    .A2(_01033_),
    .ZN(_01034_));
 NAND2_X1 _24185_ (.A1(_00958_),
    .A2(_00963_),
    .ZN(_01035_));
 NOR2_X2 _24186_ (.A1(\g_reduce0[2].adder.b[12] ),
    .A2(_00514_),
    .ZN(_01036_));
 NAND3_X2 _24187_ (.A1(_00966_),
    .A2(_00977_),
    .A3(_01036_),
    .ZN(_01037_));
 AOI21_X2 _24188_ (.A(_01037_),
    .B1(_00983_),
    .B2(_00992_),
    .ZN(_01038_));
 NOR2_X2 _24189_ (.A1(\g_reduce0[2].adder.a[12] ),
    .A2(_21412_),
    .ZN(_01039_));
 MUX2_X1 _24190_ (.A(_01039_),
    .B(_01036_),
    .S(_01004_),
    .Z(_01040_));
 AOI21_X4 _24191_ (.A(_01038_),
    .B1(_01040_),
    .B2(_01016_),
    .ZN(_01041_));
 NAND3_X4 _24192_ (.A1(_00994_),
    .A2(_01015_),
    .A3(_01039_),
    .ZN(_01042_));
 AOI21_X4 _24193_ (.A(_01035_),
    .B1(_01041_),
    .B2(_01042_),
    .ZN(_01043_));
 NOR3_X4 _24194_ (.A1(_01026_),
    .A2(_01034_),
    .A3(_01043_),
    .ZN(_01044_));
 INV_X1 _24195_ (.A(_01033_),
    .ZN(_01045_));
 INV_X1 _24196_ (.A(_00963_),
    .ZN(_01046_));
 AOI21_X4 _24197_ (.A(_01046_),
    .B1(_01041_),
    .B2(_01042_),
    .ZN(_01047_));
 AOI21_X4 _24198_ (.A(_00965_),
    .B1(_01020_),
    .B2(_01025_),
    .ZN(_01048_));
 OR4_X4 _24199_ (.A1(_00958_),
    .A2(_01045_),
    .A3(_01047_),
    .A4(_01048_),
    .ZN(_01049_));
 NAND2_X2 _24200_ (.A1(_01044_),
    .A2(_01049_),
    .ZN(_01050_));
 BUF_X4 _24201_ (.A(_21453_),
    .Z(_01051_));
 NAND2_X1 _24202_ (.A1(_00961_),
    .A2(_01051_),
    .ZN(_01052_));
 INV_X1 _24203_ (.A(_00516_),
    .ZN(_01053_));
 INV_X1 _24204_ (.A(_21421_),
    .ZN(_01054_));
 MUX2_X1 _24205_ (.A(_01053_),
    .B(_01054_),
    .S(_01018_),
    .Z(_01055_));
 INV_X1 _24206_ (.A(_00515_),
    .ZN(_01056_));
 INV_X1 _24207_ (.A(_21418_),
    .ZN(_01057_));
 MUX2_X1 _24208_ (.A(_01056_),
    .B(_01057_),
    .S(_01018_),
    .Z(_01058_));
 MUX2_X1 _24209_ (.A(_01055_),
    .B(_01058_),
    .S(_00961_),
    .Z(_01059_));
 OAI21_X1 _24210_ (.A(_01052_),
    .B1(_01059_),
    .B2(_01051_),
    .ZN(_01060_));
 INV_X1 _24211_ (.A(_01019_),
    .ZN(_01061_));
 AOI211_X2 _24212_ (.A(_00974_),
    .B(_01061_),
    .C1(_00993_),
    .C2(_00994_),
    .ZN(_01062_));
 OR3_X2 _24213_ (.A1(_21452_),
    .A2(_01023_),
    .A3(_01024_),
    .ZN(_01063_));
 OAI21_X1 _24214_ (.A(_00964_),
    .B1(_01062_),
    .B2(_01063_),
    .ZN(_01064_));
 INV_X1 _24215_ (.A(_00964_),
    .ZN(_01065_));
 NAND3_X2 _24216_ (.A1(_01065_),
    .A2(_01020_),
    .A3(_01025_),
    .ZN(_01066_));
 NAND2_X2 _24217_ (.A1(_01064_),
    .A2(_01066_),
    .ZN(_01067_));
 BUF_X1 _24218_ (.A(_01067_),
    .Z(_01068_));
 INV_X1 _24219_ (.A(_21448_),
    .ZN(_01069_));
 AOI21_X2 _24220_ (.A(_00962_),
    .B1(_01069_),
    .B2(_00997_),
    .ZN(_01070_));
 OAI221_X2 _24221_ (.A(_01005_),
    .B1(_01019_),
    .B2(_01070_),
    .C1(_01015_),
    .C2(_01016_),
    .ZN(_01071_));
 OAI21_X1 _24222_ (.A(_21417_),
    .B1(_01069_),
    .B2(_00997_),
    .ZN(_01072_));
 OAI21_X2 _24223_ (.A(_01072_),
    .B1(_00509_),
    .B2(_00952_),
    .ZN(_01073_));
 NAND2_X1 _24224_ (.A1(_00999_),
    .A2(_01073_),
    .ZN(_01074_));
 OAI22_X2 _24225_ (.A1(_00965_),
    .A2(_01071_),
    .B1(_01074_),
    .B2(_00995_),
    .ZN(_01075_));
 OR2_X1 _24226_ (.A1(\g_reduce0[2].adder.a[12] ),
    .A2(_21412_),
    .ZN(_01076_));
 INV_X1 _24227_ (.A(_01036_),
    .ZN(_01077_));
 MUX2_X1 _24228_ (.A(_01076_),
    .B(_01077_),
    .S(_01004_),
    .Z(_01078_));
 AND2_X1 _24229_ (.A1(_00992_),
    .A2(_00983_),
    .ZN(_01079_));
 OAI22_X2 _24230_ (.A1(_00994_),
    .A2(_01078_),
    .B1(_01037_),
    .B2(_01079_),
    .ZN(_01080_));
 NOR3_X1 _24231_ (.A1(_01016_),
    .A2(_00993_),
    .A3(_01076_),
    .ZN(_01081_));
 NOR3_X1 _24232_ (.A1(_00963_),
    .A2(_01080_),
    .A3(_01081_),
    .ZN(_01082_));
 NOR2_X1 _24233_ (.A1(_01019_),
    .A2(_01070_),
    .ZN(_01083_));
 AOI211_X2 _24234_ (.A(_00974_),
    .B(_01083_),
    .C1(_00993_),
    .C2(_00994_),
    .ZN(_01084_));
 AND2_X1 _24235_ (.A1(_00964_),
    .A2(_01073_),
    .ZN(_01085_));
 AOI22_X2 _24236_ (.A1(_00964_),
    .A2(_01084_),
    .B1(_01085_),
    .B2(_01017_),
    .ZN(_01086_));
 AOI211_X2 _24237_ (.A(_01047_),
    .B(_01075_),
    .C1(_01082_),
    .C2(_01086_),
    .ZN(_01087_));
 CLKBUF_X3 _24238_ (.A(_01087_),
    .Z(_01088_));
 NAND2_X1 _24239_ (.A1(_01068_),
    .A2(_01088_),
    .ZN(_01089_));
 MUX2_X1 _24240_ (.A(_00512_),
    .B(_21424_),
    .S(_01004_),
    .Z(_01090_));
 NAND2_X1 _24241_ (.A1(_01016_),
    .A2(_01090_),
    .ZN(_01091_));
 NAND3_X1 _24242_ (.A1(_21424_),
    .A2(_00994_),
    .A3(_00993_),
    .ZN(_01092_));
 NAND3_X1 _24243_ (.A1(_00512_),
    .A2(_01005_),
    .A3(_01015_),
    .ZN(_01093_));
 NAND3_X1 _24244_ (.A1(_01091_),
    .A2(_01092_),
    .A3(_01093_),
    .ZN(_01094_));
 INV_X1 _24245_ (.A(_00510_),
    .ZN(_01095_));
 AOI211_X2 _24246_ (.A(_01095_),
    .B(_00974_),
    .C1(_00993_),
    .C2(_00994_),
    .ZN(_01096_));
 INV_X1 _24247_ (.A(_21430_),
    .ZN(_01097_));
 NOR2_X1 _24248_ (.A1(_00994_),
    .A2(_01004_),
    .ZN(_01098_));
 AOI211_X2 _24249_ (.A(_01097_),
    .B(_01098_),
    .C1(_01015_),
    .C2(_00994_),
    .ZN(_01099_));
 OR2_X1 _24250_ (.A1(_01096_),
    .A2(_01099_),
    .ZN(_01100_));
 INV_X1 _24251_ (.A(_21453_),
    .ZN(_01101_));
 CLKBUF_X3 _24252_ (.A(_01101_),
    .Z(_01102_));
 MUX2_X1 _24253_ (.A(_01094_),
    .B(_01100_),
    .S(_01102_),
    .Z(_01103_));
 BUF_X4 _24254_ (.A(_01018_),
    .Z(_01104_));
 MUX2_X1 _24255_ (.A(_00513_),
    .B(_21427_),
    .S(_01104_),
    .Z(_01105_));
 NAND2_X1 _24256_ (.A1(_01051_),
    .A2(_01105_),
    .ZN(_01106_));
 AND2_X1 _24257_ (.A1(_00511_),
    .A2(_00995_),
    .ZN(_01107_));
 AOI21_X1 _24258_ (.A(_01107_),
    .B1(_01104_),
    .B2(_21433_),
    .ZN(_01108_));
 OAI21_X1 _24259_ (.A(_01106_),
    .B1(_01108_),
    .B2(_01051_),
    .ZN(_01109_));
 CLKBUF_X3 _24260_ (.A(_00960_),
    .Z(_01110_));
 MUX2_X1 _24261_ (.A(_01103_),
    .B(_01109_),
    .S(_01110_),
    .Z(_01111_));
 MUX2_X1 _24262_ (.A(_21445_),
    .B(_00505_),
    .S(_01104_),
    .Z(_01112_));
 NAND2_X1 _24263_ (.A1(_01102_),
    .A2(_01112_),
    .ZN(_01113_));
 NOR2_X1 _24264_ (.A1(_01016_),
    .A2(_01015_),
    .ZN(_01114_));
 MUX2_X1 _24265_ (.A(_00508_),
    .B(_21439_),
    .S(_01004_),
    .Z(_01115_));
 NOR2_X1 _24266_ (.A1(_01016_),
    .A2(_00993_),
    .ZN(_01116_));
 AOI222_X2 _24267_ (.A1(_21439_),
    .A2(_01114_),
    .B1(_01115_),
    .B2(_01016_),
    .C1(_01116_),
    .C2(_00508_),
    .ZN(_01117_));
 OAI21_X1 _24268_ (.A(_01113_),
    .B1(_01117_),
    .B2(_01102_),
    .ZN(_01118_));
 MUX2_X1 _24269_ (.A(_00507_),
    .B(_21436_),
    .S(_01104_),
    .Z(_01119_));
 MUX2_X1 _24270_ (.A(_00504_),
    .B(_21442_),
    .S(_01104_),
    .Z(_01120_));
 MUX2_X1 _24271_ (.A(_01119_),
    .B(_01120_),
    .S(_01102_),
    .Z(_01121_));
 MUX2_X1 _24272_ (.A(_01118_),
    .B(_01121_),
    .S(_00961_),
    .Z(_01122_));
 MUX2_X1 _24273_ (.A(_01111_),
    .B(_01122_),
    .S(_01068_),
    .Z(_01123_));
 OAI22_X1 _24274_ (.A1(_01060_),
    .A2(_01089_),
    .B1(_01123_),
    .B2(_01088_),
    .ZN(_01124_));
 NAND2_X1 _24275_ (.A1(_01050_),
    .A2(_01124_),
    .ZN(_21520_));
 INV_X1 _24276_ (.A(_21520_),
    .ZN(_21517_));
 MUX2_X1 _24277_ (.A(_00515_),
    .B(_21418_),
    .S(_01018_),
    .Z(_01125_));
 AOI21_X2 _24278_ (.A(_01051_),
    .B1(_01125_),
    .B2(_01110_),
    .ZN(_01126_));
 NAND3_X1 _24279_ (.A1(_01068_),
    .A2(_01088_),
    .A3(_01126_),
    .ZN(_01127_));
 AOI21_X4 _24280_ (.A(_01065_),
    .B1(_01020_),
    .B2(_01025_),
    .ZN(_01128_));
 NOR3_X4 _24281_ (.A1(_00964_),
    .A2(_01062_),
    .A3(_01063_),
    .ZN(_01129_));
 NOR2_X4 _24282_ (.A1(_01128_),
    .A2(_01129_),
    .ZN(_01130_));
 MUX2_X1 _24283_ (.A(_00516_),
    .B(_21421_),
    .S(_01018_),
    .Z(_01131_));
 MUX2_X1 _24284_ (.A(_01131_),
    .B(_01105_),
    .S(_01102_),
    .Z(_01132_));
 MUX2_X1 _24285_ (.A(_01103_),
    .B(_01132_),
    .S(_00961_),
    .Z(_01133_));
 NAND2_X1 _24286_ (.A1(_01130_),
    .A2(_01133_),
    .ZN(_01134_));
 MUX2_X1 _24287_ (.A(_01108_),
    .B(_01117_),
    .S(_01102_),
    .Z(_01135_));
 NOR2_X1 _24288_ (.A1(_01110_),
    .A2(_01135_),
    .ZN(_01136_));
 AOI21_X1 _24289_ (.A(_01136_),
    .B1(_01121_),
    .B2(_01110_),
    .ZN(_01137_));
 OAI21_X1 _24290_ (.A(_01134_),
    .B1(_01137_),
    .B2(_01130_),
    .ZN(_01138_));
 OAI21_X1 _24291_ (.A(_01127_),
    .B1(_01138_),
    .B2(_01088_),
    .ZN(_01139_));
 NAND2_X2 _24292_ (.A1(_01050_),
    .A2(_01139_),
    .ZN(_14094_));
 INV_X1 _24293_ (.A(_14094_),
    .ZN(_14089_));
 AOI21_X4 _24294_ (.A(_01088_),
    .B1(_01049_),
    .B2(_01044_),
    .ZN(_01140_));
 NAND3_X2 _24295_ (.A1(_01068_),
    .A2(_01126_),
    .A3(_01140_),
    .ZN(_21472_));
 INV_X1 _24296_ (.A(_21472_),
    .ZN(_21476_));
 OAI21_X1 _24297_ (.A(_00963_),
    .B1(_01080_),
    .B2(_01081_),
    .ZN(_01141_));
 NAND2_X1 _24298_ (.A1(_00964_),
    .A2(_01073_),
    .ZN(_01142_));
 OAI22_X1 _24299_ (.A1(_01065_),
    .A2(_01071_),
    .B1(_01142_),
    .B2(_00995_),
    .ZN(_01143_));
 NAND3_X1 _24300_ (.A1(_01046_),
    .A2(_01041_),
    .A3(_01042_),
    .ZN(_01144_));
 AOI21_X1 _24301_ (.A(_01084_),
    .B1(_01073_),
    .B2(_01018_),
    .ZN(_01145_));
 OAI221_X1 _24302_ (.A(_01141_),
    .B1(_01143_),
    .B2(_01144_),
    .C1(_01145_),
    .C2(_00965_),
    .ZN(_01146_));
 CLKBUF_X3 _24303_ (.A(_01146_),
    .Z(_01147_));
 NOR4_X4 _24304_ (.A1(_00958_),
    .A2(_01045_),
    .A3(_01047_),
    .A4(_01048_),
    .ZN(_01148_));
 OR3_X4 _24305_ (.A1(_01026_),
    .A2(_01034_),
    .A3(_01043_),
    .ZN(_01149_));
 OAI21_X2 _24306_ (.A(_01147_),
    .B1(_01148_),
    .B2(_01149_),
    .ZN(_01150_));
 OR3_X1 _24307_ (.A1(_01060_),
    .A2(_01130_),
    .A3(_01150_),
    .ZN(_21465_));
 INV_X1 _24308_ (.A(_21465_),
    .ZN(_21469_));
 NOR2_X2 _24309_ (.A1(_01110_),
    .A2(_01051_),
    .ZN(_01151_));
 NOR2_X4 _24310_ (.A1(_00961_),
    .A2(_01051_),
    .ZN(_01152_));
 NOR2_X1 _24311_ (.A1(_00961_),
    .A2(_01102_),
    .ZN(_01153_));
 AOI222_X2 _24312_ (.A1(_01131_),
    .A2(_01151_),
    .B1(_01152_),
    .B2(_01094_),
    .C1(_01153_),
    .C2(_01125_),
    .ZN(_01154_));
 NAND3_X1 _24313_ (.A1(_01068_),
    .A2(_01140_),
    .A3(_01154_),
    .ZN(_21500_));
 INV_X1 _24314_ (.A(_21500_),
    .ZN(_21504_));
 NAND2_X1 _24315_ (.A1(_01110_),
    .A2(_01102_),
    .ZN(_01155_));
 NOR2_X1 _24316_ (.A1(_01068_),
    .A2(_01155_),
    .ZN(_01156_));
 NAND2_X1 _24317_ (.A1(_01051_),
    .A2(_01059_),
    .ZN(_01157_));
 MUX2_X1 _24318_ (.A(_01094_),
    .B(_01105_),
    .S(_01110_),
    .Z(_01158_));
 OAI21_X1 _24319_ (.A(_01157_),
    .B1(_01158_),
    .B2(_01051_),
    .ZN(_01159_));
 AOI21_X1 _24320_ (.A(_01156_),
    .B1(_01159_),
    .B2(_01068_),
    .ZN(_01160_));
 OR2_X1 _24321_ (.A1(_01150_),
    .A2(_01160_),
    .ZN(_21479_));
 INV_X1 _24322_ (.A(_21479_),
    .ZN(_21483_));
 NAND2_X1 _24323_ (.A1(_01130_),
    .A2(_01126_),
    .ZN(_01161_));
 OAI21_X1 _24324_ (.A(_01161_),
    .B1(_01133_),
    .B2(_01130_),
    .ZN(_01162_));
 AND2_X1 _24325_ (.A1(_01140_),
    .A2(_01162_),
    .ZN(_21486_));
 INV_X1 _24326_ (.A(_21486_),
    .ZN(_21490_));
 MUX2_X1 _24327_ (.A(_01060_),
    .B(_01111_),
    .S(_01068_),
    .Z(_01163_));
 NOR2_X1 _24328_ (.A1(_01150_),
    .A2(_01163_),
    .ZN(_21493_));
 INV_X1 _24329_ (.A(_21493_),
    .ZN(_21497_));
 NOR2_X2 _24330_ (.A1(_01110_),
    .A2(_01102_),
    .ZN(_01164_));
 AOI222_X2 _24331_ (.A1(_00513_),
    .A2(_01164_),
    .B1(_01151_),
    .B2(_00511_),
    .C1(_00507_),
    .C2(_01152_),
    .ZN(_01165_));
 AOI222_X2 _24332_ (.A1(_21427_),
    .A2(_01164_),
    .B1(_01151_),
    .B2(_21433_),
    .C1(_21436_),
    .C2(_01152_),
    .ZN(_01166_));
 MUX2_X1 _24333_ (.A(_01165_),
    .B(_01166_),
    .S(_01017_),
    .Z(_01167_));
 OAI21_X1 _24334_ (.A(_01153_),
    .B1(_01099_),
    .B2(_01096_),
    .ZN(_01168_));
 AND2_X1 _24335_ (.A1(_01167_),
    .A2(_01168_),
    .ZN(_01169_));
 MUX2_X1 _24336_ (.A(_01154_),
    .B(_01169_),
    .S(_01068_),
    .Z(_01170_));
 AND2_X1 _24337_ (.A1(_01140_),
    .A2(_01170_),
    .ZN(_21510_));
 INV_X1 _24338_ (.A(_21510_),
    .ZN(_21514_));
 NAND2_X1 _24339_ (.A1(_01110_),
    .A2(_01135_),
    .ZN(_01171_));
 MUX2_X1 _24340_ (.A(_01100_),
    .B(_01119_),
    .S(_01102_),
    .Z(_01172_));
 OAI21_X1 _24341_ (.A(_01171_),
    .B1(_01172_),
    .B2(_01110_),
    .ZN(_01173_));
 MUX2_X1 _24342_ (.A(_01159_),
    .B(_01173_),
    .S(_01068_),
    .Z(_01174_));
 NOR2_X1 _24343_ (.A1(_01088_),
    .A2(_01174_),
    .ZN(_01175_));
 OAI21_X2 _24344_ (.A(_01152_),
    .B1(_01129_),
    .B2(_01128_),
    .ZN(_01176_));
 AOI21_X1 _24345_ (.A(_01175_),
    .B1(_01176_),
    .B2(_01088_),
    .ZN(_01177_));
 NAND2_X1 _24346_ (.A1(_01050_),
    .A2(_01177_),
    .ZN(_21507_));
 INV_X1 _24347_ (.A(_21507_),
    .ZN(_21461_));
 XOR2_X2 _24348_ (.A(_00947_),
    .B(_00948_),
    .Z(_01178_));
 BUF_X4 _24349_ (.A(_01178_),
    .Z(_01179_));
 BUF_X2 _24350_ (.A(_21475_),
    .Z(_01180_));
 INV_X2 _24351_ (.A(_01180_),
    .ZN(_01181_));
 INV_X1 _24352_ (.A(_21470_),
    .ZN(_01182_));
 NOR2_X1 _24353_ (.A1(_21488_),
    .A2(_21495_),
    .ZN(_01183_));
 INV_X1 _24354_ (.A(_01183_),
    .ZN(_01184_));
 BUF_X2 _24355_ (.A(_21496_),
    .Z(_01185_));
 INV_X2 _24356_ (.A(_01185_),
    .ZN(_01186_));
 BUF_X2 _24357_ (.A(_21513_),
    .Z(_01187_));
 INV_X1 _24358_ (.A(_01187_),
    .ZN(_01188_));
 INV_X1 _24359_ (.A(_21512_),
    .ZN(_01189_));
 AOI21_X2 _24360_ (.A(_01186_),
    .B1(_01188_),
    .B2(_01189_),
    .ZN(_01190_));
 NOR2_X1 _24361_ (.A1(_21463_),
    .A2(_21512_),
    .ZN(_01191_));
 AOI21_X1 _24362_ (.A(_21457_),
    .B1(_14088_),
    .B2(_21458_),
    .ZN(_01192_));
 INV_X1 _24363_ (.A(_21464_),
    .ZN(_01193_));
 OAI21_X2 _24364_ (.A(_01191_),
    .B1(_01192_),
    .B2(_01193_),
    .ZN(_01194_));
 AOI21_X4 _24365_ (.A(_01184_),
    .B1(_01190_),
    .B2(_01194_),
    .ZN(_01195_));
 CLKBUF_X3 _24366_ (.A(_21468_),
    .Z(_01196_));
 INV_X1 _24367_ (.A(_01196_),
    .ZN(_01197_));
 BUF_X2 _24368_ (.A(_21482_),
    .Z(_01198_));
 NOR2_X1 _24369_ (.A1(_21489_),
    .A2(_21488_),
    .ZN(_01199_));
 NOR3_X2 _24370_ (.A1(_01198_),
    .A2(_21503_),
    .A3(_01199_),
    .ZN(_01200_));
 NAND2_X1 _24371_ (.A1(_01197_),
    .A2(_01200_),
    .ZN(_01201_));
 INV_X2 _24372_ (.A(_21503_),
    .ZN(_01202_));
 AOI21_X1 _24373_ (.A(_21505_),
    .B1(_21484_),
    .B2(_01202_),
    .ZN(_01203_));
 OAI221_X2 _24374_ (.A(_01182_),
    .B1(_01195_),
    .B2(_01201_),
    .C1(_01203_),
    .C2(_01196_),
    .ZN(_01204_));
 AOI21_X4 _24375_ (.A(_21477_),
    .B1(_01181_),
    .B2(_01204_),
    .ZN(_01205_));
 NOR2_X2 _24376_ (.A1(_01179_),
    .A2(_01205_),
    .ZN(_01206_));
 INV_X1 _24377_ (.A(_21467_),
    .ZN(_01207_));
 OR2_X1 _24378_ (.A1(_21491_),
    .A2(_21498_),
    .ZN(_01208_));
 NOR2_X1 _24379_ (.A1(_21502_),
    .A2(_01208_),
    .ZN(_01209_));
 INV_X2 _24380_ (.A(_21481_),
    .ZN(_01210_));
 OAI21_X2 _24381_ (.A(_01209_),
    .B1(_01210_),
    .B2(_01202_),
    .ZN(_01211_));
 NOR2_X1 _24382_ (.A1(_21508_),
    .A2(_21515_),
    .ZN(_01212_));
 AOI21_X2 _24383_ (.A(_21459_),
    .B1(_14093_),
    .B2(_21460_),
    .ZN(_01213_));
 INV_X1 _24384_ (.A(_21509_),
    .ZN(_01214_));
 OAI21_X2 _24385_ (.A(_01212_),
    .B1(_01213_),
    .B2(_01214_),
    .ZN(_01215_));
 INV_X1 _24386_ (.A(_21515_),
    .ZN(_01216_));
 AOI21_X2 _24387_ (.A(_01185_),
    .B1(_01187_),
    .B2(_01216_),
    .ZN(_01217_));
 AND2_X1 _24388_ (.A1(_01215_),
    .A2(_01217_),
    .ZN(_01218_));
 INV_X2 _24389_ (.A(_21489_),
    .ZN(_01219_));
 OAI21_X2 _24390_ (.A(_01198_),
    .B1(_21491_),
    .B2(_01219_),
    .ZN(_01220_));
 AOI21_X4 _24391_ (.A(_01202_),
    .B1(_01210_),
    .B2(_01220_),
    .ZN(_01221_));
 OAI221_X2 _24392_ (.A(_01196_),
    .B1(_01211_),
    .B2(_01218_),
    .C1(_01221_),
    .C2(_21502_),
    .ZN(_01222_));
 AOI21_X2 _24393_ (.A(_01181_),
    .B1(_01207_),
    .B2(_01222_),
    .ZN(_01223_));
 OAI21_X4 _24394_ (.A(_01179_),
    .B1(_01223_),
    .B2(_21474_),
    .ZN(_01224_));
 AOI211_X2 _24395_ (.A(_01087_),
    .B(_01176_),
    .C1(_01044_),
    .C2(_01049_),
    .ZN(_01225_));
 BUF_X4 _24396_ (.A(_01225_),
    .Z(_01226_));
 AOI21_X4 _24397_ (.A(_01206_),
    .B1(_01224_),
    .B2(_01226_),
    .ZN(_01227_));
 BUF_X4 _24398_ (.A(_01227_),
    .Z(_01228_));
 AOI21_X1 _24399_ (.A(_01180_),
    .B1(_21474_),
    .B2(_01178_),
    .ZN(_01229_));
 AOI21_X2 _24400_ (.A(_21463_),
    .B1(_14091_),
    .B2(_21464_),
    .ZN(_01230_));
 NAND2_X1 _24401_ (.A1(_01185_),
    .A2(_01187_),
    .ZN(_01231_));
 OAI221_X2 _24402_ (.A(_01183_),
    .B1(_01230_),
    .B2(_01231_),
    .C1(_01189_),
    .C2(_01186_),
    .ZN(_01232_));
 AOI221_X2 _24403_ (.A(_21505_),
    .B1(_21484_),
    .B2(_01202_),
    .C1(_01200_),
    .C2(_01232_),
    .ZN(_01233_));
 OAI21_X1 _24404_ (.A(_01182_),
    .B1(_01233_),
    .B2(_01196_),
    .ZN(_01234_));
 OAI21_X2 _24405_ (.A(_01229_),
    .B1(_01234_),
    .B2(_01179_),
    .ZN(_01235_));
 XNOR2_X2 _24406_ (.A(_00947_),
    .B(_00948_),
    .ZN(_01236_));
 BUF_X4 _24407_ (.A(_01236_),
    .Z(_01237_));
 BUF_X4 _24408_ (.A(_01237_),
    .Z(_01238_));
 NAND2_X2 _24409_ (.A1(_21477_),
    .A2(_01238_),
    .ZN(_01239_));
 NOR3_X1 _24410_ (.A1(_21474_),
    .A2(_21467_),
    .A3(_01238_),
    .ZN(_01240_));
 AOI21_X2 _24411_ (.A(_21508_),
    .B1(_14095_),
    .B2(_21509_),
    .ZN(_01241_));
 OAI21_X1 _24412_ (.A(_01216_),
    .B1(_01241_),
    .B2(_01187_),
    .ZN(_01242_));
 AND2_X1 _24413_ (.A1(_01186_),
    .A2(_01242_),
    .ZN(_01243_));
 OAI22_X2 _24414_ (.A1(_21502_),
    .A2(_01221_),
    .B1(_01243_),
    .B2(_01211_),
    .ZN(_01244_));
 OAI21_X2 _24415_ (.A(_01240_),
    .B1(_01244_),
    .B2(_01197_),
    .ZN(_01245_));
 AND3_X1 _24416_ (.A1(_01235_),
    .A2(_01239_),
    .A3(_01245_),
    .ZN(_01246_));
 XNOR2_X2 _24417_ (.A(_01226_),
    .B(_01246_),
    .ZN(_01247_));
 NAND2_X1 _24418_ (.A1(_01237_),
    .A2(_01233_),
    .ZN(_01248_));
 OAI221_X2 _24419_ (.A(_01178_),
    .B1(_01211_),
    .B2(_01243_),
    .C1(_01221_),
    .C2(_21502_),
    .ZN(_01249_));
 AND3_X2 _24420_ (.A1(_01196_),
    .A2(_01248_),
    .A3(_01249_),
    .ZN(_01250_));
 AOI21_X4 _24421_ (.A(_01196_),
    .B1(_01248_),
    .B2(_01249_),
    .ZN(_01251_));
 OR2_X4 _24422_ (.A1(_01250_),
    .A2(_01251_),
    .ZN(_01252_));
 INV_X1 _24423_ (.A(_21498_),
    .ZN(_01253_));
 OR2_X1 _24424_ (.A1(_01185_),
    .A2(_01187_),
    .ZN(_01254_));
 OAI221_X2 _24425_ (.A(_01253_),
    .B1(_01241_),
    .B2(_01254_),
    .C1(_01216_),
    .C2(_01185_),
    .ZN(_01255_));
 AOI211_X2 _24426_ (.A(_21491_),
    .B(_01236_),
    .C1(_01255_),
    .C2(_01219_),
    .ZN(_01256_));
 OR2_X1 _24427_ (.A1(_21489_),
    .A2(_21488_),
    .ZN(_01257_));
 AND3_X1 _24428_ (.A1(_01237_),
    .A2(_01257_),
    .A3(_01232_),
    .ZN(_01258_));
 OR3_X2 _24429_ (.A1(_01198_),
    .A2(_01256_),
    .A3(_01258_),
    .ZN(_01259_));
 OAI21_X2 _24430_ (.A(_01198_),
    .B1(_01256_),
    .B2(_01258_),
    .ZN(_01260_));
 OAI21_X1 _24431_ (.A(_01189_),
    .B1(_01230_),
    .B2(_01188_),
    .ZN(_01261_));
 AND2_X1 _24432_ (.A1(_01237_),
    .A2(_01261_),
    .ZN(_01262_));
 NOR2_X2 _24433_ (.A1(_01237_),
    .A2(_01242_),
    .ZN(_01263_));
 OR3_X2 _24434_ (.A1(_01186_),
    .A2(_01262_),
    .A3(_01263_),
    .ZN(_01264_));
 OAI21_X4 _24435_ (.A(_01186_),
    .B1(_01262_),
    .B2(_01263_),
    .ZN(_01265_));
 NAND4_X4 _24436_ (.A1(_01259_),
    .A2(_01260_),
    .A3(_01264_),
    .A4(_01265_),
    .ZN(_01266_));
 NOR2_X4 _24437_ (.A1(_01252_),
    .A2(_01266_),
    .ZN(_01267_));
 OAI21_X2 _24438_ (.A(_01202_),
    .B1(_01210_),
    .B2(_01237_),
    .ZN(_01268_));
 OR2_X1 _24439_ (.A1(_01198_),
    .A2(_01199_),
    .ZN(_01269_));
 OAI21_X1 _24440_ (.A(_21503_),
    .B1(_01195_),
    .B2(_01269_),
    .ZN(_01270_));
 AOI21_X1 _24441_ (.A(_01208_),
    .B1(_01215_),
    .B2(_01217_),
    .ZN(_01271_));
 OR2_X1 _24442_ (.A1(_01236_),
    .A2(_01220_),
    .ZN(_01272_));
 OAI22_X2 _24443_ (.A1(_21484_),
    .A2(_01178_),
    .B1(_01271_),
    .B2(_01272_),
    .ZN(_01273_));
 MUX2_X2 _24444_ (.A(_01268_),
    .B(_01270_),
    .S(_01273_),
    .Z(_01274_));
 NOR3_X2 _24445_ (.A1(_01195_),
    .A2(_01269_),
    .A3(_01268_),
    .ZN(_01275_));
 NOR3_X2 _24446_ (.A1(_01202_),
    .A2(_01210_),
    .A3(_01237_),
    .ZN(_01276_));
 NOR2_X4 _24447_ (.A1(_01275_),
    .A2(_01276_),
    .ZN(_01277_));
 AOI21_X2 _24448_ (.A(_21498_),
    .B1(_01215_),
    .B2(_01217_),
    .ZN(_01278_));
 OR2_X1 _24449_ (.A1(_21495_),
    .A2(_01178_),
    .ZN(_01279_));
 AND2_X1 _24450_ (.A1(_01194_),
    .A2(_01190_),
    .ZN(_01280_));
 OAI22_X4 _24451_ (.A1(_01237_),
    .A2(_01278_),
    .B1(_01279_),
    .B2(_01280_),
    .ZN(_01281_));
 XNOR2_X2 _24452_ (.A(_21489_),
    .B(_01281_),
    .ZN(_01282_));
 AND2_X2 _24453_ (.A1(_01259_),
    .A2(_01260_),
    .ZN(_01283_));
 AOI22_X4 _24454_ (.A1(_01274_),
    .A2(_01277_),
    .B1(_01282_),
    .B2(_01283_),
    .ZN(_01284_));
 AND2_X1 _24455_ (.A1(_01238_),
    .A2(_01204_),
    .ZN(_01285_));
 AND3_X2 _24456_ (.A1(_01207_),
    .A2(_01179_),
    .A3(_01222_),
    .ZN(_01286_));
 NOR3_X4 _24457_ (.A1(_01181_),
    .A2(_01285_),
    .A3(_01286_),
    .ZN(_01287_));
 NAND2_X2 _24458_ (.A1(_01238_),
    .A2(_01204_),
    .ZN(_01288_));
 NAND3_X2 _24459_ (.A1(_01207_),
    .A2(_01179_),
    .A3(_01222_),
    .ZN(_01289_));
 AOI21_X4 _24460_ (.A(_01180_),
    .B1(_01288_),
    .B2(_01289_),
    .ZN(_01290_));
 OAI22_X4 _24461_ (.A1(_01252_),
    .A2(_01284_),
    .B1(_01287_),
    .B2(_01290_),
    .ZN(_01291_));
 OAI21_X4 _24462_ (.A(_01247_),
    .B1(_01267_),
    .B2(_01291_),
    .ZN(_01292_));
 XOR2_X2 _24463_ (.A(_14091_),
    .B(_21464_),
    .Z(_01293_));
 NAND2_X1 _24464_ (.A1(_01237_),
    .A2(_01293_),
    .ZN(_01294_));
 XOR2_X2 _24465_ (.A(_14095_),
    .B(_21509_),
    .Z(_01295_));
 NAND2_X1 _24466_ (.A1(_01178_),
    .A2(_01295_),
    .ZN(_01296_));
 NAND2_X2 _24467_ (.A1(_01294_),
    .A2(_01296_),
    .ZN(_01297_));
 MUX2_X2 _24468_ (.A(_21519_),
    .B(_21521_),
    .S(_01178_),
    .Z(_01298_));
 NOR2_X1 _24469_ (.A1(_01297_),
    .A2(_01298_),
    .ZN(_01299_));
 NAND2_X2 _24470_ (.A1(_01179_),
    .A2(_01299_),
    .ZN(_01300_));
 NAND2_X1 _24471_ (.A1(_00961_),
    .A2(_01101_),
    .ZN(_01301_));
 AND3_X1 _24472_ (.A1(_01091_),
    .A2(_01092_),
    .A3(_01093_),
    .ZN(_01302_));
 NAND2_X1 _24473_ (.A1(_00960_),
    .A2(_01051_),
    .ZN(_01303_));
 OAI222_X2 _24474_ (.A1(_01055_),
    .A2(_01301_),
    .B1(_01155_),
    .B2(_01302_),
    .C1(_01303_),
    .C2(_01058_),
    .ZN(_01304_));
 NOR3_X4 _24475_ (.A1(_01130_),
    .A2(_01147_),
    .A3(_01304_),
    .ZN(_01305_));
 AOI211_X4 _24476_ (.A(_01128_),
    .B(_01129_),
    .C1(_01167_),
    .C2(_01168_),
    .ZN(_01306_));
 OAI22_X1 _24477_ (.A1(_00505_),
    .A2(_01301_),
    .B1(_01303_),
    .B2(_21442_),
    .ZN(_01307_));
 OAI22_X1 _24478_ (.A1(_21445_),
    .A2(_01301_),
    .B1(_01303_),
    .B2(_00504_),
    .ZN(_01308_));
 MUX2_X1 _24479_ (.A(_01307_),
    .B(_01308_),
    .S(_00995_),
    .Z(_01309_));
 AOI221_X4 _24480_ (.A(_01309_),
    .B1(_01066_),
    .B2(_01064_),
    .C1(_01164_),
    .C2(_01117_),
    .ZN(_01310_));
 NOR3_X4 _24481_ (.A1(_01087_),
    .A2(_01306_),
    .A3(_01310_),
    .ZN(_01311_));
 NOR3_X4 _24482_ (.A1(_01300_),
    .A2(_01305_),
    .A3(_01311_),
    .ZN(_01312_));
 NOR3_X2 _24483_ (.A1(_01179_),
    .A2(_01293_),
    .A3(_01298_),
    .ZN(_01313_));
 OAI221_X2 _24484_ (.A(_01313_),
    .B1(_01129_),
    .B2(_01128_),
    .C1(_01149_),
    .C2(_01148_),
    .ZN(_01314_));
 AOI21_X1 _24485_ (.A(_01309_),
    .B1(_01117_),
    .B2(_01164_),
    .ZN(_01315_));
 MUX2_X1 _24486_ (.A(_01304_),
    .B(_01315_),
    .S(_01147_),
    .Z(_01316_));
 NOR2_X2 _24487_ (.A1(_01314_),
    .A2(_01316_),
    .ZN(_01317_));
 INV_X1 _24488_ (.A(_21508_),
    .ZN(_01318_));
 OAI21_X2 _24489_ (.A(_01318_),
    .B1(_01214_),
    .B2(_01213_),
    .ZN(_01319_));
 NOR2_X1 _24490_ (.A1(_21463_),
    .A2(_01178_),
    .ZN(_01320_));
 OR2_X1 _24491_ (.A1(_01193_),
    .A2(_01192_),
    .ZN(_01321_));
 AOI22_X4 _24492_ (.A1(_01178_),
    .A2(_01319_),
    .B1(_01320_),
    .B2(_01321_),
    .ZN(_01322_));
 XNOR2_X2 _24493_ (.A(_01188_),
    .B(_01322_),
    .ZN(_01323_));
 AND2_X1 _24494_ (.A1(_14092_),
    .A2(_01237_),
    .ZN(_01324_));
 AOI21_X4 _24495_ (.A(_01324_),
    .B1(_01178_),
    .B2(_14096_),
    .ZN(_01325_));
 AND2_X2 _24496_ (.A1(_01294_),
    .A2(_01296_),
    .ZN(_01326_));
 AOI21_X4 _24497_ (.A(_01323_),
    .B1(_01325_),
    .B2(_01326_),
    .ZN(_01327_));
 NAND3_X1 _24498_ (.A1(_01130_),
    .A2(_01169_),
    .A3(_01313_),
    .ZN(_01328_));
 OAI221_X2 _24499_ (.A(_01327_),
    .B1(_01328_),
    .B2(_01150_),
    .C1(_01050_),
    .C2(_01300_),
    .ZN(_01329_));
 NOR4_X4 _24500_ (.A1(_01291_),
    .A2(_01312_),
    .A3(_01317_),
    .A4(_01329_),
    .ZN(_01330_));
 OAI21_X4 _24501_ (.A(_01228_),
    .B1(_01292_),
    .B2(_01330_),
    .ZN(_21523_));
 INV_X1 _24502_ (.A(_21523_),
    .ZN(_21525_));
 BUF_X2 _24503_ (.A(_21528_),
    .Z(_01331_));
 OR2_X1 _24504_ (.A1(_01206_),
    .A2(_01246_),
    .ZN(_01332_));
 NOR2_X4 _24505_ (.A1(_01250_),
    .A2(_01251_),
    .ZN(_01333_));
 NAND3_X1 _24506_ (.A1(_01181_),
    .A2(_01288_),
    .A3(_01289_),
    .ZN(_01334_));
 OAI21_X1 _24507_ (.A(_01180_),
    .B1(_01285_),
    .B2(_01286_),
    .ZN(_01335_));
 NAND2_X2 _24508_ (.A1(_01259_),
    .A2(_01260_),
    .ZN(_01336_));
 AOI21_X4 _24509_ (.A(_01336_),
    .B1(_01274_),
    .B2(_01277_),
    .ZN(_01337_));
 AND4_X2 _24510_ (.A1(_01333_),
    .A2(_01334_),
    .A3(_01335_),
    .A4(_01337_),
    .ZN(_01338_));
 AND2_X2 _24511_ (.A1(_01264_),
    .A2(_01265_),
    .ZN(_01339_));
 XNOR2_X2 _24512_ (.A(_01219_),
    .B(_01281_),
    .ZN(_01340_));
 XNOR2_X2 _24513_ (.A(_01187_),
    .B(_01322_),
    .ZN(_01341_));
 NAND4_X4 _24514_ (.A1(_01339_),
    .A2(_01340_),
    .A3(_01326_),
    .A4(_01341_),
    .ZN(_01342_));
 AOI21_X1 _24515_ (.A(_01332_),
    .B1(_01338_),
    .B2(_01342_),
    .ZN(_01343_));
 NAND3_X4 _24516_ (.A1(_01235_),
    .A2(_01239_),
    .A3(_01245_),
    .ZN(_01344_));
 OR2_X1 _24517_ (.A1(_01224_),
    .A2(_01344_),
    .ZN(_01345_));
 AOI21_X1 _24518_ (.A(_01345_),
    .B1(_01338_),
    .B2(_01342_),
    .ZN(_01346_));
 MUX2_X2 _24519_ (.A(_01343_),
    .B(_01346_),
    .S(_01225_),
    .Z(_01347_));
 XNOR2_X2 _24520_ (.A(_01331_),
    .B(_01347_),
    .ZN(_01348_));
 INV_X2 _24521_ (.A(_01348_),
    .ZN(_01349_));
 BUF_X8 _24522_ (.A(_01349_),
    .Z(_01350_));
 CLKBUF_X3 _24523_ (.A(_01350_),
    .Z(_21549_));
 INV_X1 _24524_ (.A(_01332_),
    .ZN(_01351_));
 INV_X1 _24525_ (.A(_01345_),
    .ZN(_01352_));
 MUX2_X2 _24526_ (.A(_01351_),
    .B(_01352_),
    .S(_01226_),
    .Z(_01353_));
 CLKBUF_X3 _24527_ (.A(_01353_),
    .Z(_01354_));
 BUF_X1 _24528_ (.A(_21524_),
    .Z(_01355_));
 NOR2_X1 _24529_ (.A1(_01355_),
    .A2(_01298_),
    .ZN(_01356_));
 OAI22_X1 _24530_ (.A1(_01331_),
    .A2(_01338_),
    .B1(_01354_),
    .B2(_01356_),
    .ZN(_01357_));
 INV_X1 _24531_ (.A(_01331_),
    .ZN(_01358_));
 NAND2_X2 _24532_ (.A1(_01342_),
    .A2(_01338_),
    .ZN(_01359_));
 NOR2_X1 _24533_ (.A1(_01358_),
    .A2(_01359_),
    .ZN(_01360_));
 NAND3_X2 _24534_ (.A1(_01180_),
    .A2(_01288_),
    .A3(_01289_),
    .ZN(_01361_));
 OAI21_X2 _24535_ (.A(_01181_),
    .B1(_01285_),
    .B2(_01286_),
    .ZN(_01362_));
 AND2_X1 _24536_ (.A1(_21519_),
    .A2(_01238_),
    .ZN(_01363_));
 AOI21_X4 _24537_ (.A(_01363_),
    .B1(_01179_),
    .B2(_21521_),
    .ZN(_01364_));
 MUX2_X1 _24538_ (.A(_14096_),
    .B(_14092_),
    .S(_01238_),
    .Z(_01365_));
 CLKBUF_X3 _24539_ (.A(_01365_),
    .Z(_01366_));
 NAND2_X1 _24540_ (.A1(_01364_),
    .A2(_01366_),
    .ZN(_01367_));
 NAND3_X1 _24541_ (.A1(_01326_),
    .A2(_01341_),
    .A3(_01367_),
    .ZN(_01368_));
 NAND3_X1 _24542_ (.A1(_01339_),
    .A2(_01340_),
    .A3(_01368_),
    .ZN(_01369_));
 AOI221_X2 _24543_ (.A(_01252_),
    .B1(_01361_),
    .B2(_01362_),
    .C1(_01337_),
    .C2(_01369_),
    .ZN(_01370_));
 NOR2_X2 _24544_ (.A1(_01252_),
    .A2(_01284_),
    .ZN(_01371_));
 NOR4_X1 _24545_ (.A1(_01250_),
    .A2(_01251_),
    .A3(_01266_),
    .A4(_01327_),
    .ZN(_01372_));
 OR2_X1 _24546_ (.A1(_01371_),
    .A2(_01372_),
    .ZN(_01373_));
 OR3_X1 _24547_ (.A1(_01250_),
    .A2(_01251_),
    .A3(_01266_),
    .ZN(_01374_));
 CLKBUF_X3 _24548_ (.A(_01374_),
    .Z(_01375_));
 NAND2_X1 _24549_ (.A1(_01238_),
    .A2(_01299_),
    .ZN(_01376_));
 NOR4_X1 _24550_ (.A1(_01087_),
    .A2(_01375_),
    .A3(_01310_),
    .A4(_01376_),
    .ZN(_01377_));
 AOI21_X1 _24551_ (.A(_01306_),
    .B1(_01049_),
    .B2(_01044_),
    .ZN(_01378_));
 AOI221_X2 _24552_ (.A(_01376_),
    .B1(_01066_),
    .B2(_01064_),
    .C1(_01044_),
    .C2(_01049_),
    .ZN(_01379_));
 NOR3_X1 _24553_ (.A1(_01147_),
    .A2(_01304_),
    .A3(_01375_),
    .ZN(_01380_));
 AOI221_X2 _24554_ (.A(_01373_),
    .B1(_01377_),
    .B2(_01378_),
    .C1(_01379_),
    .C2(_01380_),
    .ZN(_01381_));
 NOR3_X2 _24555_ (.A1(_01238_),
    .A2(_01295_),
    .A3(_01298_),
    .ZN(_01382_));
 NAND2_X2 _24556_ (.A1(_01267_),
    .A2(_01382_),
    .ZN(_01383_));
 NOR2_X4 _24557_ (.A1(_01149_),
    .A2(_01148_),
    .ZN(_01384_));
 NAND3_X2 _24558_ (.A1(_01067_),
    .A2(_01088_),
    .A3(_01154_),
    .ZN(_01385_));
 OR3_X2 _24559_ (.A1(_01087_),
    .A2(_01306_),
    .A3(_01310_),
    .ZN(_01386_));
 AOI21_X4 _24560_ (.A(_01384_),
    .B1(_01385_),
    .B2(_01386_),
    .ZN(_01387_));
 OAI211_X4 _24561_ (.A(_01370_),
    .B(_01381_),
    .C1(_01383_),
    .C2(_01387_),
    .ZN(_01388_));
 AOI21_X1 _24562_ (.A(_01357_),
    .B1(_01360_),
    .B2(_01388_),
    .ZN(_01389_));
 MUX2_X2 _24563_ (.A(_01332_),
    .B(_01345_),
    .S(_01226_),
    .Z(_01390_));
 OAI21_X1 _24564_ (.A(_01267_),
    .B1(_01312_),
    .B2(_01317_),
    .ZN(_01391_));
 AOI21_X1 _24565_ (.A(_01291_),
    .B1(_01329_),
    .B2(_01267_),
    .ZN(_01392_));
 AOI21_X1 _24566_ (.A(_01147_),
    .B1(_01154_),
    .B2(_01067_),
    .ZN(_01393_));
 OAI21_X2 _24567_ (.A(_01179_),
    .B1(_01306_),
    .B2(_01393_),
    .ZN(_01394_));
 OAI221_X2 _24568_ (.A(_01238_),
    .B1(_01305_),
    .B2(_01311_),
    .C1(_01148_),
    .C2(_01149_),
    .ZN(_01395_));
 AOI22_X1 _24569_ (.A1(_01044_),
    .A2(_01049_),
    .B1(_01147_),
    .B2(_01310_),
    .ZN(_01396_));
 OR2_X2 _24570_ (.A1(_01238_),
    .A2(_01396_),
    .ZN(_01397_));
 NAND3_X4 _24571_ (.A1(_01394_),
    .A2(_01395_),
    .A3(_01397_),
    .ZN(_01398_));
 BUF_X4 _24572_ (.A(_14098_),
    .Z(_01399_));
 AOI221_X2 _24573_ (.A(_01390_),
    .B1(_01391_),
    .B2(_01392_),
    .C1(_01398_),
    .C2(_01399_),
    .ZN(_01400_));
 AOI21_X1 _24574_ (.A(_01356_),
    .B1(_01366_),
    .B2(_01355_),
    .ZN(_01401_));
 NOR2_X1 _24575_ (.A1(_01354_),
    .A2(_01401_),
    .ZN(_01402_));
 CLKBUF_X3 _24576_ (.A(_01399_),
    .Z(_01403_));
 NAND3_X1 _24577_ (.A1(_01403_),
    .A2(_01364_),
    .A3(_01354_),
    .ZN(_01404_));
 OR4_X1 _24578_ (.A1(_01291_),
    .A2(_01312_),
    .A3(_01317_),
    .A4(_01329_),
    .ZN(_01405_));
 CLKBUF_X3 _24579_ (.A(_01405_),
    .Z(_01406_));
 XNOR2_X2 _24580_ (.A(_01226_),
    .B(_01344_),
    .ZN(_01407_));
 NOR2_X4 _24581_ (.A1(_01287_),
    .A2(_01290_),
    .ZN(_01408_));
 NOR2_X2 _24582_ (.A1(_01371_),
    .A2(_01408_),
    .ZN(_01409_));
 AOI21_X2 _24583_ (.A(_01407_),
    .B1(_01375_),
    .B2(_01409_),
    .ZN(_01410_));
 BUF_X4 _24584_ (.A(_01410_),
    .Z(_01411_));
 AOI21_X1 _24585_ (.A(_01404_),
    .B1(_01406_),
    .B2(_01411_),
    .ZN(_01412_));
 NOR4_X2 _24586_ (.A1(_01389_),
    .A2(_01400_),
    .A3(_01402_),
    .A4(_01412_),
    .ZN(_01413_));
 INV_X1 _24587_ (.A(_01355_),
    .ZN(_01414_));
 CLKBUF_X3 _24588_ (.A(_01414_),
    .Z(_01415_));
 NOR2_X1 _24589_ (.A1(_01415_),
    .A2(_01298_),
    .ZN(_01416_));
 NOR2_X1 _24590_ (.A1(_01354_),
    .A2(_01416_),
    .ZN(_01417_));
 CLKBUF_X3 _24591_ (.A(_01355_),
    .Z(_01418_));
 OAI21_X1 _24592_ (.A(_01417_),
    .B1(_01398_),
    .B2(_01418_),
    .ZN(_01419_));
 NAND2_X2 _24593_ (.A1(_01361_),
    .A2(_01362_),
    .ZN(_01420_));
 NAND3_X2 _24594_ (.A1(_01333_),
    .A2(_01420_),
    .A3(_01337_),
    .ZN(_01421_));
 AND2_X1 _24595_ (.A1(_01342_),
    .A2(_01353_),
    .ZN(_01422_));
 AOI22_X4 _24596_ (.A1(_01421_),
    .A2(_01353_),
    .B1(_01388_),
    .B2(_01422_),
    .ZN(_01423_));
 OAI222_X2 _24597_ (.A1(_01252_),
    .A2(_01284_),
    .B1(_01287_),
    .B2(_01290_),
    .C1(_01327_),
    .C2(_01375_),
    .ZN(_01424_));
 NAND2_X1 _24598_ (.A1(_01344_),
    .A2(_01424_),
    .ZN(_01425_));
 NAND2_X1 _24599_ (.A1(_01246_),
    .A2(_01424_),
    .ZN(_01426_));
 MUX2_X2 _24600_ (.A(_01425_),
    .B(_01426_),
    .S(_01226_),
    .Z(_01427_));
 NAND4_X2 _24601_ (.A1(_01394_),
    .A2(_01395_),
    .A3(_01397_),
    .A4(_01427_),
    .ZN(_01428_));
 INV_X2 _24602_ (.A(_01399_),
    .ZN(_01429_));
 NAND4_X2 _24603_ (.A1(_01067_),
    .A2(_01147_),
    .A3(_01152_),
    .A4(_01224_),
    .ZN(_01430_));
 OAI22_X4 _24604_ (.A1(_01179_),
    .A2(_01205_),
    .B1(_01430_),
    .B2(_01384_),
    .ZN(_01431_));
 NOR2_X2 _24605_ (.A1(_01429_),
    .A2(_01431_),
    .ZN(_01432_));
 XNOR2_X1 _24606_ (.A(_01331_),
    .B(_01359_),
    .ZN(_01433_));
 BUF_X4 _24607_ (.A(_01390_),
    .Z(_01434_));
 AOI21_X1 _24608_ (.A(_01433_),
    .B1(_01416_),
    .B2(_01434_),
    .ZN(_01435_));
 NAND3_X1 _24609_ (.A1(_01428_),
    .A2(_01432_),
    .A3(_01435_),
    .ZN(_01436_));
 OAI21_X1 _24610_ (.A(_01419_),
    .B1(_01423_),
    .B2(_01436_),
    .ZN(_01437_));
 NAND2_X1 _24611_ (.A1(_01413_),
    .A2(_01437_),
    .ZN(_01438_));
 INV_X1 _24612_ (.A(_01438_),
    .ZN(_21531_));
 NOR2_X1 _24613_ (.A1(_00951_),
    .A2(_00957_),
    .ZN(_01439_));
 AOI22_X2 _24614_ (.A1(\g_reduce0[2].adder.b[0] ),
    .A2(_00951_),
    .B1(_01439_),
    .B2(\g_reduce0[2].adder.a[0] ),
    .ZN(_01440_));
 INV_X2 _24615_ (.A(_00950_),
    .ZN(_01441_));
 CLKBUF_X3 _24616_ (.A(_01441_),
    .Z(_01442_));
 NAND2_X1 _24617_ (.A1(_01442_),
    .A2(_00957_),
    .ZN(_01443_));
 NAND2_X2 _24618_ (.A1(_01418_),
    .A2(_01434_),
    .ZN(_01444_));
 CLKBUF_X3 _24619_ (.A(_01407_),
    .Z(_01445_));
 NAND2_X2 _24620_ (.A1(_01338_),
    .A2(_01353_),
    .ZN(_01446_));
 INV_X1 _24621_ (.A(_01359_),
    .ZN(_01447_));
 AOI21_X2 _24622_ (.A(_01446_),
    .B1(_01388_),
    .B2(_01447_),
    .ZN(_01448_));
 OAI21_X1 _24623_ (.A(_01432_),
    .B1(_01398_),
    .B2(_01350_),
    .ZN(_01449_));
 NAND3_X1 _24624_ (.A1(_01411_),
    .A2(_01297_),
    .A3(_01406_),
    .ZN(_01450_));
 OAI21_X1 _24625_ (.A(_01323_),
    .B1(_01330_),
    .B2(_01292_),
    .ZN(_01451_));
 AND2_X1 _24626_ (.A1(_01450_),
    .A2(_01451_),
    .ZN(_01452_));
 AOI21_X1 _24627_ (.A(_01449_),
    .B1(_01452_),
    .B2(_21549_),
    .ZN(_01453_));
 CLKBUF_X3 _24628_ (.A(_01429_),
    .Z(_01454_));
 NOR2_X1 _24629_ (.A1(_01292_),
    .A2(_01330_),
    .ZN(_01455_));
 CLKBUF_X3 _24630_ (.A(_01348_),
    .Z(_01456_));
 NAND2_X1 _24631_ (.A1(_01455_),
    .A2(_01456_),
    .ZN(_01457_));
 MUX2_X1 _24632_ (.A(_01366_),
    .B(_01364_),
    .S(_01455_),
    .Z(_01458_));
 NAND2_X1 _24633_ (.A1(_01454_),
    .A2(_21549_),
    .ZN(_01459_));
 OAI22_X1 _24634_ (.A1(_01454_),
    .A2(_01457_),
    .B1(_01458_),
    .B2(_01459_),
    .ZN(_01460_));
 OAI21_X1 _24635_ (.A(_01448_),
    .B1(_01453_),
    .B2(_01460_),
    .ZN(_01461_));
 AOI21_X1 _24636_ (.A(_01431_),
    .B1(_01247_),
    .B2(_01333_),
    .ZN(_01462_));
 AOI21_X2 _24637_ (.A(_01348_),
    .B1(_01462_),
    .B2(_01408_),
    .ZN(_01463_));
 NAND2_X2 _24638_ (.A1(_01264_),
    .A2(_01265_),
    .ZN(_01464_));
 AND2_X1 _24639_ (.A1(_01344_),
    .A2(_01291_),
    .ZN(_01465_));
 AND2_X1 _24640_ (.A1(_01246_),
    .A2(_01291_),
    .ZN(_01466_));
 MUX2_X2 _24641_ (.A(_01465_),
    .B(_01466_),
    .S(_01226_),
    .Z(_01467_));
 MUX2_X1 _24642_ (.A(_01282_),
    .B(_01464_),
    .S(_01467_),
    .Z(_01468_));
 NOR2_X1 _24643_ (.A1(_21549_),
    .A2(_01468_),
    .ZN(_01469_));
 NOR3_X1 _24644_ (.A1(_01403_),
    .A2(_01463_),
    .A3(_01469_),
    .ZN(_01470_));
 NOR2_X1 _24645_ (.A1(_01333_),
    .A2(_01408_),
    .ZN(_01471_));
 NOR3_X1 _24646_ (.A1(_01226_),
    .A2(_01246_),
    .A3(_01471_),
    .ZN(_01472_));
 NOR4_X1 _24647_ (.A1(_01150_),
    .A2(_01176_),
    .A3(_01344_),
    .A4(_01471_),
    .ZN(_01473_));
 NAND2_X1 _24648_ (.A1(_01274_),
    .A2(_01277_),
    .ZN(_01474_));
 OAI33_X1 _24649_ (.A1(_01407_),
    .A2(_01283_),
    .A3(_01409_),
    .B1(_01472_),
    .B2(_01473_),
    .B3(_01474_),
    .ZN(_01475_));
 AND2_X1 _24650_ (.A1(_01456_),
    .A2(_01475_),
    .ZN(_01476_));
 AOI21_X1 _24651_ (.A(_01470_),
    .B1(_01476_),
    .B2(_01403_),
    .ZN(_01477_));
 AOI21_X2 _24652_ (.A(_01445_),
    .B1(_01461_),
    .B2(_01477_),
    .ZN(_01478_));
 BUF_X4 _24653_ (.A(_01431_),
    .Z(_01479_));
 OAI21_X4 _24654_ (.A(_01444_),
    .B1(_01478_),
    .B2(_01479_),
    .ZN(_01480_));
 NOR2_X1 _24655_ (.A1(_01479_),
    .A2(_01359_),
    .ZN(_01481_));
 AOI22_X4 _24656_ (.A1(_01228_),
    .A2(_01446_),
    .B1(_01481_),
    .B2(_01388_),
    .ZN(_01482_));
 INV_X1 _24657_ (.A(_01482_),
    .ZN(_21553_));
 MUX2_X1 _24658_ (.A(_01336_),
    .B(_01282_),
    .S(_01467_),
    .Z(_01483_));
 NOR2_X1 _24659_ (.A1(_01454_),
    .A2(_01483_),
    .ZN(_01484_));
 NAND2_X1 _24660_ (.A1(_01341_),
    .A2(_01467_),
    .ZN(_01485_));
 AOI221_X2 _24661_ (.A(_01399_),
    .B1(_01410_),
    .B2(_01323_),
    .C1(_01485_),
    .C2(_01464_),
    .ZN(_01486_));
 NOR3_X1 _24662_ (.A1(_21549_),
    .A2(_01484_),
    .A3(_01486_),
    .ZN(_01487_));
 NAND3_X1 _24663_ (.A1(_01454_),
    .A2(_01474_),
    .A3(_01408_),
    .ZN(_01488_));
 NAND2_X1 _24664_ (.A1(_01403_),
    .A2(_01420_),
    .ZN(_01489_));
 AOI21_X1 _24665_ (.A(_01445_),
    .B1(_01488_),
    .B2(_01489_),
    .ZN(_01490_));
 NOR4_X1 _24666_ (.A1(_01403_),
    .A2(_01479_),
    .A3(_01247_),
    .A4(_01252_),
    .ZN(_01491_));
 AOI221_X2 _24667_ (.A(_01403_),
    .B1(_01228_),
    .B2(_01252_),
    .C1(_01274_),
    .C2(_01277_),
    .ZN(_01492_));
 NOR4_X1 _24668_ (.A1(_01456_),
    .A2(_01490_),
    .A3(_01491_),
    .A4(_01492_),
    .ZN(_01493_));
 NOR2_X1 _24669_ (.A1(_01415_),
    .A2(_01445_),
    .ZN(_01494_));
 NOR2_X1 _24670_ (.A1(_01418_),
    .A2(_01479_),
    .ZN(_01495_));
 OAI221_X1 _24671_ (.A(_21553_),
    .B1(_01487_),
    .B2(_01493_),
    .C1(_01494_),
    .C2(_01495_),
    .ZN(_01496_));
 NAND2_X1 _24672_ (.A1(_21526_),
    .A2(_01456_),
    .ZN(_01497_));
 NOR2_X1 _24673_ (.A1(_01399_),
    .A2(_01431_),
    .ZN(_01498_));
 NAND2_X1 _24674_ (.A1(_01350_),
    .A2(_01498_),
    .ZN(_01499_));
 NAND3_X1 _24675_ (.A1(_01228_),
    .A2(_01445_),
    .A3(_01364_),
    .ZN(_01500_));
 AND2_X1 _24676_ (.A1(_01227_),
    .A2(_01427_),
    .ZN(_01501_));
 NAND3_X1 _24677_ (.A1(_01227_),
    .A2(_01409_),
    .A3(_01364_),
    .ZN(_01502_));
 NOR2_X2 _24678_ (.A1(_01375_),
    .A2(_01300_),
    .ZN(_01503_));
 NAND3_X1 _24679_ (.A1(_01385_),
    .A2(_01386_),
    .A3(_01503_),
    .ZN(_01504_));
 OR3_X1 _24680_ (.A1(_01375_),
    .A2(_01314_),
    .A3(_01316_),
    .ZN(_01505_));
 OAI21_X1 _24681_ (.A(_01341_),
    .B1(_01366_),
    .B2(_01297_),
    .ZN(_01506_));
 AND3_X1 _24682_ (.A1(_01130_),
    .A2(_01169_),
    .A3(_01313_),
    .ZN(_01507_));
 AOI221_X2 _24683_ (.A(_01506_),
    .B1(_01507_),
    .B2(_01140_),
    .C1(_01384_),
    .C2(_01382_),
    .ZN(_01508_));
 OAI211_X2 _24684_ (.A(_01504_),
    .B(_01505_),
    .C1(_01375_),
    .C2(_01508_),
    .ZN(_01509_));
 OAI221_X2 _24685_ (.A(_01500_),
    .B1(_01501_),
    .B2(_01398_),
    .C1(_01502_),
    .C2(_01509_),
    .ZN(_01510_));
 NAND2_X1 _24686_ (.A1(_01350_),
    .A2(_01432_),
    .ZN(_01511_));
 NAND4_X1 _24687_ (.A1(_01226_),
    .A2(_01246_),
    .A3(_01408_),
    .A4(_01325_),
    .ZN(_01512_));
 NAND3_X1 _24688_ (.A1(_01344_),
    .A2(_01408_),
    .A3(_01325_),
    .ZN(_01513_));
 OAI221_X2 _24689_ (.A(_01512_),
    .B1(_01366_),
    .B2(_01227_),
    .C1(_01226_),
    .C2(_01513_),
    .ZN(_01514_));
 NOR2_X1 _24690_ (.A1(_01479_),
    .A2(_01326_),
    .ZN(_01515_));
 OAI21_X2 _24691_ (.A(_01381_),
    .B1(_01383_),
    .B2(_01387_),
    .ZN(_01516_));
 NOR2_X1 _24692_ (.A1(_01445_),
    .A2(_01366_),
    .ZN(_01517_));
 AOI221_X2 _24693_ (.A(_01514_),
    .B1(_01515_),
    .B2(_01427_),
    .C1(_01516_),
    .C2(_01517_),
    .ZN(_01518_));
 OAI221_X2 _24694_ (.A(_01497_),
    .B1(_01499_),
    .B2(_01510_),
    .C1(_01511_),
    .C2(_01518_),
    .ZN(_01519_));
 NAND3_X1 _24695_ (.A1(_01482_),
    .A2(_01519_),
    .A3(_01494_),
    .ZN(_01520_));
 NOR2_X1 _24696_ (.A1(_01415_),
    .A2(_01228_),
    .ZN(_01521_));
 AND2_X1 _24697_ (.A1(_01482_),
    .A2(_01495_),
    .ZN(_01522_));
 AOI221_X1 _24698_ (.A(_01521_),
    .B1(_01522_),
    .B2(_01519_),
    .C1(_01415_),
    .C2(_01445_),
    .ZN(_01523_));
 AND3_X1 _24699_ (.A1(_01496_),
    .A2(_01520_),
    .A3(_01523_),
    .ZN(_01524_));
 MUX2_X1 _24700_ (.A(_01333_),
    .B(_01420_),
    .S(_01355_),
    .Z(_01525_));
 NOR2_X1 _24701_ (.A1(_01354_),
    .A2(_01525_),
    .ZN(_01526_));
 NAND2_X1 _24702_ (.A1(_01358_),
    .A2(_01347_),
    .ZN(_01527_));
 NAND2_X1 _24703_ (.A1(_01337_),
    .A2(_01369_),
    .ZN(_01528_));
 NAND3_X1 _24704_ (.A1(_01333_),
    .A2(_01420_),
    .A3(_01528_),
    .ZN(_01529_));
 NOR2_X1 _24705_ (.A1(_01359_),
    .A2(_01529_),
    .ZN(_01530_));
 OAI21_X1 _24706_ (.A(_01331_),
    .B1(_01434_),
    .B2(_01530_),
    .ZN(_01531_));
 OAI21_X1 _24707_ (.A(_01527_),
    .B1(_01531_),
    .B2(_21523_),
    .ZN(_01532_));
 NAND4_X2 _24708_ (.A1(_01399_),
    .A2(_01411_),
    .A3(_01406_),
    .A4(_01398_),
    .ZN(_01533_));
 OAI22_X2 _24709_ (.A1(_01454_),
    .A2(_01298_),
    .B1(_01330_),
    .B2(_01292_),
    .ZN(_01534_));
 AOI21_X1 _24710_ (.A(_01446_),
    .B1(_01533_),
    .B2(_01534_),
    .ZN(_01535_));
 AOI21_X1 _24711_ (.A(_01333_),
    .B1(_01408_),
    .B2(_01247_),
    .ZN(_01536_));
 OAI21_X1 _24712_ (.A(_01403_),
    .B1(_01445_),
    .B2(_01474_),
    .ZN(_01537_));
 OAI221_X1 _24713_ (.A(_21549_),
    .B1(_01536_),
    .B2(_01537_),
    .C1(_01483_),
    .C2(_01403_),
    .ZN(_01538_));
 NOR2_X1 _24714_ (.A1(_01399_),
    .A2(_01366_),
    .ZN(_01539_));
 NOR2_X1 _24715_ (.A1(_01429_),
    .A2(_01341_),
    .ZN(_01540_));
 OAI21_X1 _24716_ (.A(_01408_),
    .B1(_01539_),
    .B2(_01540_),
    .ZN(_01541_));
 INV_X1 _24717_ (.A(_01541_),
    .ZN(_01542_));
 MUX2_X1 _24718_ (.A(_01464_),
    .B(_01297_),
    .S(_01429_),
    .Z(_01543_));
 MUX2_X1 _24719_ (.A(_01542_),
    .B(_01543_),
    .S(_01445_),
    .Z(_01544_));
 AOI21_X2 _24720_ (.A(_01429_),
    .B1(_01464_),
    .B2(_01409_),
    .ZN(_01545_));
 OAI21_X1 _24721_ (.A(_01323_),
    .B1(_01371_),
    .B2(_01267_),
    .ZN(_01546_));
 OAI21_X1 _24722_ (.A(_01545_),
    .B1(_01546_),
    .B2(_01445_),
    .ZN(_01547_));
 OAI21_X1 _24723_ (.A(_01429_),
    .B1(_01326_),
    .B2(_01424_),
    .ZN(_01548_));
 AOI211_X2 _24724_ (.A(_01407_),
    .B(_01366_),
    .C1(_01546_),
    .C2(_01545_),
    .ZN(_01549_));
 AOI221_X2 _24725_ (.A(_01544_),
    .B1(_01547_),
    .B2(_01548_),
    .C1(_01549_),
    .C2(_01516_),
    .ZN(_01550_));
 OAI21_X1 _24726_ (.A(_01538_),
    .B1(_01550_),
    .B2(_21549_),
    .ZN(_01551_));
 NOR2_X1 _24727_ (.A1(_01273_),
    .A2(_01268_),
    .ZN(_01552_));
 OR2_X1 _24728_ (.A1(_01195_),
    .A2(_01269_),
    .ZN(_01553_));
 AND3_X1 _24729_ (.A1(_21503_),
    .A2(_01553_),
    .A3(_01273_),
    .ZN(_01554_));
 OR2_X1 _24730_ (.A1(_01275_),
    .A2(_01276_),
    .ZN(_01555_));
 NOR2_X1 _24731_ (.A1(_01219_),
    .A2(_01281_),
    .ZN(_01556_));
 AND2_X1 _24732_ (.A1(_01219_),
    .A2(_01281_),
    .ZN(_01557_));
 OAI33_X1 _24733_ (.A1(_01552_),
    .A2(_01554_),
    .A3(_01555_),
    .B1(_01556_),
    .B2(_01557_),
    .B3(_01336_),
    .ZN(_01558_));
 AOI21_X1 _24734_ (.A(_01372_),
    .B1(_01558_),
    .B2(_01333_),
    .ZN(_01559_));
 AND2_X1 _24735_ (.A1(_01370_),
    .A2(_01559_),
    .ZN(_01560_));
 OR4_X1 _24736_ (.A1(_01088_),
    .A2(_01375_),
    .A3(_01310_),
    .A4(_01376_),
    .ZN(_01561_));
 OAI22_X2 _24737_ (.A1(_01149_),
    .A2(_01148_),
    .B1(_01067_),
    .B2(_01169_),
    .ZN(_01562_));
 NAND3_X1 _24738_ (.A1(_01088_),
    .A2(_01154_),
    .A3(_01267_),
    .ZN(_01563_));
 OAI221_X2 _24739_ (.A(_01560_),
    .B1(_01561_),
    .B2(_01562_),
    .C1(_01314_),
    .C2(_01563_),
    .ZN(_01564_));
 OAI21_X2 _24740_ (.A(_01050_),
    .B1(_01305_),
    .B2(_01311_),
    .ZN(_01565_));
 AOI21_X4 _24741_ (.A(_01564_),
    .B1(_01503_),
    .B2(_01565_),
    .ZN(_01566_));
 NAND2_X1 _24742_ (.A1(_01342_),
    .A2(_01353_),
    .ZN(_01567_));
 OAI22_X4 _24743_ (.A1(_01338_),
    .A2(_01390_),
    .B1(_01566_),
    .B2(_01567_),
    .ZN(_01568_));
 AOI221_X2 _24744_ (.A(_01526_),
    .B1(_01532_),
    .B2(_01535_),
    .C1(_01551_),
    .C2(_01568_),
    .ZN(_01569_));
 AOI21_X1 _24745_ (.A(_01445_),
    .B1(_01479_),
    .B2(_01415_),
    .ZN(_01570_));
 AOI21_X1 _24746_ (.A(_01570_),
    .B1(_01420_),
    .B2(_01415_),
    .ZN(_01571_));
 OAI211_X2 _24747_ (.A(_01323_),
    .B(_01456_),
    .C1(_01330_),
    .C2(_01292_),
    .ZN(_01572_));
 NAND4_X1 _24748_ (.A1(_01411_),
    .A2(_01297_),
    .A3(_01406_),
    .A4(_01456_),
    .ZN(_01573_));
 NAND3_X1 _24749_ (.A1(_01228_),
    .A2(_01350_),
    .A3(_01475_),
    .ZN(_01574_));
 NAND4_X1 _24750_ (.A1(_01454_),
    .A2(_01572_),
    .A3(_01573_),
    .A4(_01574_),
    .ZN(_01575_));
 NAND2_X1 _24751_ (.A1(_01475_),
    .A2(_01498_),
    .ZN(_01576_));
 OAI21_X1 _24752_ (.A(_01228_),
    .B1(_01468_),
    .B2(_01454_),
    .ZN(_01577_));
 AOI221_X2 _24753_ (.A(_01423_),
    .B1(_01463_),
    .B2(_01576_),
    .C1(_01577_),
    .C2(_01456_),
    .ZN(_01578_));
 NOR2_X1 _24754_ (.A1(_01479_),
    .A2(_01364_),
    .ZN(_01579_));
 NAND4_X1 _24755_ (.A1(_01411_),
    .A2(_01406_),
    .A3(_01350_),
    .A4(_01579_),
    .ZN(_01580_));
 OAI21_X1 _24756_ (.A(_01325_),
    .B1(_01330_),
    .B2(_01292_),
    .ZN(_01581_));
 AND4_X1 _24757_ (.A1(_01394_),
    .A2(_01395_),
    .A3(_01397_),
    .A4(_01427_),
    .ZN(_01582_));
 OAI221_X2 _24758_ (.A(_01580_),
    .B1(_01511_),
    .B2(_01581_),
    .C1(_01582_),
    .C2(_01499_),
    .ZN(_01583_));
 AOI221_X2 _24759_ (.A(_01571_),
    .B1(_01575_),
    .B2(_01578_),
    .C1(_01583_),
    .C2(_01448_),
    .ZN(_01584_));
 OR2_X1 _24760_ (.A1(_01569_),
    .A2(_01584_),
    .ZN(_01585_));
 NOR2_X1 _24761_ (.A1(_01524_),
    .A2(_01585_),
    .ZN(_01586_));
 NAND2_X1 _24762_ (.A1(_21526_),
    .A2(_01350_),
    .ZN(_01587_));
 NAND2_X1 _24763_ (.A1(_01354_),
    .A2(_01350_),
    .ZN(_01588_));
 OAI33_X1 _24764_ (.A1(_01434_),
    .A2(_21553_),
    .A3(_01587_),
    .B1(_01588_),
    .B2(_01484_),
    .B3(_01486_),
    .ZN(_01589_));
 NAND2_X1 _24765_ (.A1(_01399_),
    .A2(_01227_),
    .ZN(_01590_));
 NAND2_X1 _24766_ (.A1(_01454_),
    .A2(_01228_),
    .ZN(_01591_));
 OAI22_X2 _24767_ (.A1(_01590_),
    .A2(_01518_),
    .B1(_01510_),
    .B2(_01591_),
    .ZN(_01592_));
 NOR2_X1 _24768_ (.A1(_21549_),
    .A2(_01423_),
    .ZN(_01593_));
 NOR2_X1 _24769_ (.A1(_01418_),
    .A2(_01336_),
    .ZN(_01594_));
 AOI21_X1 _24770_ (.A(_01594_),
    .B1(_01474_),
    .B2(_01418_),
    .ZN(_01595_));
 AOI221_X2 _24771_ (.A(_01589_),
    .B1(_01592_),
    .B2(_01593_),
    .C1(_01434_),
    .C2(_01595_),
    .ZN(_01596_));
 BUF_X1 _24772_ (.A(_01354_),
    .Z(_01597_));
 MUX2_X1 _24773_ (.A(_01333_),
    .B(_01474_),
    .S(_01414_),
    .Z(_01598_));
 NOR2_X1 _24774_ (.A1(_01597_),
    .A2(_01598_),
    .ZN(_01599_));
 AOI22_X1 _24775_ (.A1(_01432_),
    .A2(_01475_),
    .B1(_01498_),
    .B2(_01468_),
    .ZN(_01600_));
 NOR2_X1 _24776_ (.A1(_01421_),
    .A2(_01434_),
    .ZN(_01601_));
 OAI21_X1 _24777_ (.A(_01601_),
    .B1(_01566_),
    .B2(_01359_),
    .ZN(_01602_));
 NAND2_X1 _24778_ (.A1(_01428_),
    .A2(_01432_),
    .ZN(_01603_));
 OAI21_X1 _24779_ (.A(_01600_),
    .B1(_01602_),
    .B2(_01603_),
    .ZN(_01604_));
 NOR2_X1 _24780_ (.A1(_01434_),
    .A2(_01456_),
    .ZN(_01605_));
 OAI22_X1 _24781_ (.A1(_01292_),
    .A2(_01330_),
    .B1(_01539_),
    .B2(_01540_),
    .ZN(_01606_));
 NAND4_X1 _24782_ (.A1(_01454_),
    .A2(_01411_),
    .A3(_01298_),
    .A4(_01406_),
    .ZN(_01607_));
 NAND4_X1 _24783_ (.A1(_01403_),
    .A2(_01411_),
    .A3(_01297_),
    .A4(_01406_),
    .ZN(_01608_));
 NAND3_X1 _24784_ (.A1(_01606_),
    .A2(_01607_),
    .A3(_01608_),
    .ZN(_01609_));
 AOI221_X2 _24785_ (.A(_01599_),
    .B1(_01604_),
    .B2(_01605_),
    .C1(_01593_),
    .C2(_01609_),
    .ZN(_01610_));
 NOR2_X1 _24786_ (.A1(_01596_),
    .A2(_01610_),
    .ZN(_01611_));
 AOI21_X1 _24787_ (.A(_01354_),
    .B1(_01366_),
    .B2(_01415_),
    .ZN(_01612_));
 OR2_X1 _24788_ (.A1(_01568_),
    .A2(_01612_),
    .ZN(_01613_));
 OAI221_X2 _24789_ (.A(_01613_),
    .B1(_01612_),
    .B2(_01583_),
    .C1(_01297_),
    .C2(_01444_),
    .ZN(_01614_));
 OAI21_X1 _24790_ (.A(_01434_),
    .B1(_01297_),
    .B2(_01418_),
    .ZN(_01615_));
 NOR2_X1 _24791_ (.A1(_01415_),
    .A2(_01354_),
    .ZN(_01616_));
 AOI21_X2 _24792_ (.A(_01615_),
    .B1(_01616_),
    .B2(_01341_),
    .ZN(_01617_));
 AOI21_X4 _24793_ (.A(_01617_),
    .B1(_01519_),
    .B2(_01568_),
    .ZN(_01618_));
 MUX2_X1 _24794_ (.A(_01339_),
    .B(_01341_),
    .S(_01414_),
    .Z(_01619_));
 NOR2_X1 _24795_ (.A1(_01354_),
    .A2(_01619_),
    .ZN(_01620_));
 NOR3_X1 _24796_ (.A1(_01399_),
    .A2(_01479_),
    .A3(_01364_),
    .ZN(_01621_));
 NAND4_X1 _24797_ (.A1(_01411_),
    .A2(_01406_),
    .A3(_01349_),
    .A4(_01621_),
    .ZN(_01622_));
 NAND4_X1 _24798_ (.A1(_01411_),
    .A2(_01406_),
    .A3(_01348_),
    .A4(_01432_),
    .ZN(_01623_));
 NAND3_X1 _24799_ (.A1(_01228_),
    .A2(_01350_),
    .A3(_01539_),
    .ZN(_01624_));
 OAI211_X2 _24800_ (.A(_01622_),
    .B(_01623_),
    .C1(_01455_),
    .C2(_01624_),
    .ZN(_01625_));
 NOR2_X1 _24801_ (.A1(_01423_),
    .A2(_01449_),
    .ZN(_01626_));
 NAND3_X1 _24802_ (.A1(_21549_),
    .A2(_01450_),
    .A3(_01451_),
    .ZN(_01627_));
 AOI221_X2 _24803_ (.A(_01620_),
    .B1(_01625_),
    .B2(_01568_),
    .C1(_01626_),
    .C2(_01627_),
    .ZN(_01628_));
 NOR4_X2 _24804_ (.A1(_01438_),
    .A2(_01614_),
    .A3(_01618_),
    .A4(_01628_),
    .ZN(_01629_));
 NOR4_X1 _24805_ (.A1(_01479_),
    .A2(_01456_),
    .A3(_01423_),
    .A4(_01550_),
    .ZN(_01630_));
 AOI21_X1 _24806_ (.A(_01597_),
    .B1(_01339_),
    .B2(_01415_),
    .ZN(_01631_));
 AOI211_X2 _24807_ (.A(_01350_),
    .B(_01423_),
    .C1(_01533_),
    .C2(_01534_),
    .ZN(_01632_));
 OR3_X1 _24808_ (.A1(_01630_),
    .A2(_01631_),
    .A3(_01632_),
    .ZN(_01633_));
 OAI21_X1 _24809_ (.A(_01616_),
    .B1(_01340_),
    .B2(_01283_),
    .ZN(_01634_));
 NAND2_X1 _24810_ (.A1(_01414_),
    .A2(_01340_),
    .ZN(_01635_));
 AOI211_X2 _24811_ (.A(_01331_),
    .B(_01347_),
    .C1(_01635_),
    .C2(_01390_),
    .ZN(_01636_));
 AND2_X1 _24812_ (.A1(_01331_),
    .A2(_01347_),
    .ZN(_01637_));
 OAI22_X1 _24813_ (.A1(_01582_),
    .A2(_01591_),
    .B1(_01636_),
    .B2(_01637_),
    .ZN(_01638_));
 NAND3_X1 _24814_ (.A1(_01399_),
    .A2(_01228_),
    .A3(_01325_),
    .ZN(_01639_));
 AOI21_X1 _24815_ (.A(_01639_),
    .B1(_01406_),
    .B2(_01411_),
    .ZN(_01640_));
 NOR4_X1 _24816_ (.A1(_01292_),
    .A2(_01364_),
    .A3(_01330_),
    .A4(_01590_),
    .ZN(_01641_));
 NOR3_X1 _24817_ (.A1(_01638_),
    .A2(_01640_),
    .A3(_01641_),
    .ZN(_01642_));
 MUX2_X1 _24818_ (.A(_01340_),
    .B(_01339_),
    .S(_01467_),
    .Z(_01643_));
 AOI21_X1 _24819_ (.A(_01479_),
    .B1(_01643_),
    .B2(_01403_),
    .ZN(_01644_));
 OAI21_X1 _24820_ (.A(_01568_),
    .B1(_01644_),
    .B2(_01456_),
    .ZN(_01645_));
 NAND2_X1 _24821_ (.A1(_01434_),
    .A2(_01635_),
    .ZN(_01646_));
 AND3_X1 _24822_ (.A1(_01454_),
    .A2(_21549_),
    .A3(_01646_),
    .ZN(_01647_));
 AOI221_X2 _24823_ (.A(_01642_),
    .B1(_01645_),
    .B2(_01646_),
    .C1(_01452_),
    .C2(_01647_),
    .ZN(_01648_));
 AND3_X1 _24824_ (.A1(_01633_),
    .A2(_01634_),
    .A3(_01648_),
    .ZN(_01649_));
 AND3_X1 _24825_ (.A1(_01611_),
    .A2(_01629_),
    .A3(_01649_),
    .ZN(_01650_));
 NAND2_X1 _24826_ (.A1(_01586_),
    .A2(_01650_),
    .ZN(_01651_));
 XOR2_X2 _24827_ (.A(_01480_),
    .B(_01651_),
    .Z(_01652_));
 BUF_X4 _24828_ (.A(_01652_),
    .Z(_21536_));
 OAI21_X1 _24829_ (.A(_01597_),
    .B1(_01482_),
    .B2(_01587_),
    .ZN(_01653_));
 NAND2_X1 _24830_ (.A1(_01437_),
    .A2(_01653_),
    .ZN(_01654_));
 MUX2_X1 _24831_ (.A(_01654_),
    .B(_01437_),
    .S(_01413_),
    .Z(_01655_));
 NOR2_X1 _24832_ (.A1(_21536_),
    .A2(_01655_),
    .ZN(_01656_));
 AOI21_X1 _24833_ (.A(_01656_),
    .B1(_21536_),
    .B2(_21533_),
    .ZN(_01657_));
 OAI21_X2 _24834_ (.A(_01440_),
    .B1(_01443_),
    .B2(_01657_),
    .ZN(_00064_));
 NOR2_X1 _24835_ (.A1(\g_reduce0[2].adder.b[1] ),
    .A2(_01442_),
    .ZN(_01658_));
 NAND2_X1 _24836_ (.A1(_21533_),
    .A2(_00957_),
    .ZN(_01659_));
 XNOR2_X1 _24837_ (.A(_21532_),
    .B(_01618_),
    .ZN(_01660_));
 NAND2_X1 _24838_ (.A1(_00957_),
    .A2(_01660_),
    .ZN(_01661_));
 MUX2_X1 _24839_ (.A(_01659_),
    .B(_01661_),
    .S(_21536_),
    .Z(_01662_));
 NOR4_X4 _24840_ (.A1(_00952_),
    .A2(\g_reduce0[2].adder.b[12] ),
    .A3(_00953_),
    .A4(_00954_),
    .ZN(_01663_));
 AOI21_X1 _24841_ (.A(_00951_),
    .B1(_01663_),
    .B2(\g_reduce0[2].adder.a[1] ),
    .ZN(_01664_));
 AOI21_X2 _24842_ (.A(_01658_),
    .B1(_01662_),
    .B2(_01664_),
    .ZN(_00071_));
 NOR2_X1 _24843_ (.A1(\g_reduce0[2].adder.b[2] ),
    .A2(_01442_),
    .ZN(_01665_));
 OR3_X1 _24844_ (.A1(_01438_),
    .A2(_01614_),
    .A3(_01618_),
    .ZN(_01666_));
 XOR2_X2 _24845_ (.A(_01666_),
    .B(_01628_),
    .Z(_01667_));
 NAND2_X1 _24846_ (.A1(_00957_),
    .A2(_01667_),
    .ZN(_01668_));
 MUX2_X1 _24847_ (.A(_01661_),
    .B(_01668_),
    .S(_21536_),
    .Z(_01669_));
 AOI21_X1 _24848_ (.A(_00951_),
    .B1(_01663_),
    .B2(\g_reduce0[2].adder.a[2] ),
    .ZN(_01670_));
 AOI21_X2 _24849_ (.A(_01665_),
    .B1(_01669_),
    .B2(_01670_),
    .ZN(_00072_));
 INV_X1 _24850_ (.A(_21532_),
    .ZN(_01671_));
 NOR3_X2 _24851_ (.A1(_01671_),
    .A2(_01618_),
    .A3(_01628_),
    .ZN(_01672_));
 OAI21_X1 _24852_ (.A(_01633_),
    .B1(_01444_),
    .B2(_01282_),
    .ZN(_01673_));
 XNOR2_X1 _24853_ (.A(_01672_),
    .B(_01673_),
    .ZN(_01674_));
 MUX2_X1 _24854_ (.A(_01667_),
    .B(_01674_),
    .S(_21536_),
    .Z(_01675_));
 MUX2_X1 _24855_ (.A(\g_reduce0[2].adder.a[3] ),
    .B(_01675_),
    .S(_00957_),
    .Z(_01676_));
 MUX2_X1 _24856_ (.A(\g_reduce0[2].adder.b[3] ),
    .B(_01676_),
    .S(_01442_),
    .Z(_00073_));
 NOR3_X1 _24857_ (.A1(_01666_),
    .A2(_01628_),
    .A3(_01673_),
    .ZN(_01677_));
 INV_X1 _24858_ (.A(_01648_),
    .ZN(_01678_));
 AOI21_X1 _24859_ (.A(_01678_),
    .B1(_01616_),
    .B2(_01283_),
    .ZN(_01679_));
 XOR2_X1 _24860_ (.A(_01677_),
    .B(_01679_),
    .Z(_01680_));
 MUX2_X1 _24861_ (.A(_01674_),
    .B(_01680_),
    .S(_21536_),
    .Z(_01681_));
 MUX2_X1 _24862_ (.A(\g_reduce0[2].adder.a[4] ),
    .B(_01681_),
    .S(_00956_),
    .Z(_01682_));
 MUX2_X1 _24863_ (.A(\g_reduce0[2].adder.b[4] ),
    .B(_01682_),
    .S(_01442_),
    .Z(_00074_));
 NAND2_X1 _24864_ (.A1(_01649_),
    .A2(_01672_),
    .ZN(_01683_));
 XOR2_X2 _24865_ (.A(_01596_),
    .B(_01683_),
    .Z(_01684_));
 MUX2_X1 _24866_ (.A(_01680_),
    .B(_01684_),
    .S(_01652_),
    .Z(_01685_));
 MUX2_X1 _24867_ (.A(\g_reduce0[2].adder.a[5] ),
    .B(_01685_),
    .S(_00956_),
    .Z(_01686_));
 MUX2_X1 _24868_ (.A(\g_reduce0[2].adder.b[5] ),
    .B(_01686_),
    .S(_01442_),
    .Z(_00075_));
 NAND2_X1 _24869_ (.A1(\g_reduce0[2].adder.b[6] ),
    .A2(_00951_),
    .ZN(_01687_));
 OAI21_X1 _24870_ (.A(_01442_),
    .B1(_00957_),
    .B2(\g_reduce0[2].adder.a[6] ),
    .ZN(_01688_));
 NAND3_X2 _24871_ (.A1(_01611_),
    .A2(_01629_),
    .A3(_01649_),
    .ZN(_01689_));
 NAND2_X1 _24872_ (.A1(_01629_),
    .A2(_01649_),
    .ZN(_01690_));
 OAI21_X1 _24873_ (.A(_01610_),
    .B1(_01690_),
    .B2(_01596_),
    .ZN(_01691_));
 NAND2_X1 _24874_ (.A1(_01689_),
    .A2(_01691_),
    .ZN(_01692_));
 OAI21_X1 _24875_ (.A(_00957_),
    .B1(_01480_),
    .B2(_01692_),
    .ZN(_01693_));
 INV_X1 _24876_ (.A(_21536_),
    .ZN(_01694_));
 AOI21_X1 _24877_ (.A(_01693_),
    .B1(_01684_),
    .B2(_01694_),
    .ZN(_01695_));
 OAI21_X2 _24878_ (.A(_01687_),
    .B1(_01688_),
    .B2(_01695_),
    .ZN(_00076_));
 NOR2_X1 _24879_ (.A1(\g_reduce0[2].adder.b[7] ),
    .A2(_01442_),
    .ZN(_01696_));
 AOI21_X1 _24880_ (.A(_00951_),
    .B1(_01663_),
    .B2(\g_reduce0[2].adder.a[7] ),
    .ZN(_01697_));
 OAI21_X1 _24881_ (.A(_01691_),
    .B1(_01689_),
    .B2(_01586_),
    .ZN(_01698_));
 NAND2_X1 _24882_ (.A1(_01480_),
    .A2(_01698_),
    .ZN(_01699_));
 NAND3_X1 _24883_ (.A1(_01611_),
    .A2(_01649_),
    .A3(_01672_),
    .ZN(_01700_));
 XNOR2_X1 _24884_ (.A(_01569_),
    .B(_01700_),
    .ZN(_01701_));
 NAND2_X1 _24885_ (.A1(_21536_),
    .A2(_01701_),
    .ZN(_01702_));
 NOR3_X1 _24886_ (.A1(_01480_),
    .A2(_01524_),
    .A3(_01585_),
    .ZN(_01703_));
 NAND2_X1 _24887_ (.A1(_01650_),
    .A2(_01703_),
    .ZN(_01704_));
 NAND4_X1 _24888_ (.A1(_00957_),
    .A2(_01699_),
    .A3(_01702_),
    .A4(_01704_),
    .ZN(_01705_));
 AOI21_X1 _24889_ (.A(_01696_),
    .B1(_01697_),
    .B2(_01705_),
    .ZN(_00077_));
 NOR2_X1 _24890_ (.A1(\g_reduce0[2].adder.b[8] ),
    .A2(_01442_),
    .ZN(_01706_));
 AOI21_X1 _24891_ (.A(_00951_),
    .B1(_01663_),
    .B2(\g_reduce0[2].adder.a[8] ),
    .ZN(_01707_));
 XNOR2_X1 _24892_ (.A(_01480_),
    .B(_01524_),
    .ZN(_01708_));
 AOI211_X2 _24893_ (.A(_01585_),
    .B(_01689_),
    .C1(_01683_),
    .C2(_01708_),
    .ZN(_01709_));
 NAND2_X1 _24894_ (.A1(_01480_),
    .A2(_01701_),
    .ZN(_01710_));
 OAI21_X1 _24895_ (.A(_01584_),
    .B1(_01689_),
    .B2(_01569_),
    .ZN(_01711_));
 OAI21_X1 _24896_ (.A(_01710_),
    .B1(_01711_),
    .B2(_01480_),
    .ZN(_01712_));
 OR3_X1 _24897_ (.A1(_01663_),
    .A2(_01709_),
    .A3(_01712_),
    .ZN(_01713_));
 AOI21_X2 _24898_ (.A(_01706_),
    .B1(_01707_),
    .B2(_01713_),
    .ZN(_00078_));
 NOR2_X1 _24899_ (.A1(\g_reduce0[2].adder.b[9] ),
    .A2(_01442_),
    .ZN(_01714_));
 AOI21_X1 _24900_ (.A(_00951_),
    .B1(_01663_),
    .B2(\g_reduce0[2].adder.a[9] ),
    .ZN(_01715_));
 NOR2_X1 _24901_ (.A1(_01585_),
    .A2(_01700_),
    .ZN(_01716_));
 XNOR2_X1 _24902_ (.A(_01524_),
    .B(_01716_),
    .ZN(_01717_));
 NOR2_X1 _24903_ (.A1(_01569_),
    .A2(_01689_),
    .ZN(_01718_));
 XNOR2_X1 _24904_ (.A(_01584_),
    .B(_01718_),
    .ZN(_01719_));
 AOI22_X1 _24905_ (.A1(_21536_),
    .A2(_01717_),
    .B1(_01719_),
    .B2(_01480_),
    .ZN(_01720_));
 OR2_X1 _24906_ (.A1(_01663_),
    .A2(_01720_),
    .ZN(_01721_));
 AOI21_X2 _24907_ (.A(_01714_),
    .B1(_01715_),
    .B2(_01721_),
    .ZN(_00079_));
 INV_X1 _24908_ (.A(_21534_),
    .ZN(_21540_));
 MUX2_X1 _24909_ (.A(\g_reduce0[2].adder.a[10] ),
    .B(_21539_),
    .S(_00956_),
    .Z(_01722_));
 MUX2_X2 _24910_ (.A(\g_reduce0[2].adder.b[10] ),
    .B(_01722_),
    .S(_01441_),
    .Z(_00065_));
 MUX2_X1 _24911_ (.A(\g_reduce0[2].adder.a[11] ),
    .B(_21547_),
    .S(_00956_),
    .Z(_01723_));
 MUX2_X2 _24912_ (.A(_00952_),
    .B(_01723_),
    .S(_01441_),
    .Z(_00066_));
 MUX2_X2 _24913_ (.A(_21412_),
    .B(_00514_),
    .S(_01018_),
    .Z(_01724_));
 NAND2_X1 _24914_ (.A1(_01418_),
    .A2(_21541_),
    .ZN(_01725_));
 XOR2_X1 _24915_ (.A(_01724_),
    .B(_01725_),
    .Z(_01726_));
 XOR2_X1 _24916_ (.A(_14100_),
    .B(_21551_),
    .Z(_01727_));
 MUX2_X1 _24917_ (.A(_01726_),
    .B(_01727_),
    .S(_01597_),
    .Z(_01728_));
 XOR2_X1 _24918_ (.A(_21546_),
    .B(_01728_),
    .Z(_01729_));
 MUX2_X1 _24919_ (.A(\g_reduce0[2].adder.a[12] ),
    .B(_01729_),
    .S(_00956_),
    .Z(_01730_));
 MUX2_X2 _24920_ (.A(\g_reduce0[2].adder.b[12] ),
    .B(_01730_),
    .S(_01441_),
    .Z(_00067_));
 INV_X1 _24921_ (.A(_14102_),
    .ZN(_14099_));
 MUX2_X1 _24922_ (.A(_21409_),
    .B(_00517_),
    .S(_01018_),
    .Z(_01731_));
 MUX2_X1 _24923_ (.A(_21415_),
    .B(_00509_),
    .S(_01018_),
    .Z(_01732_));
 NOR4_X1 _24924_ (.A1(_01415_),
    .A2(_21534_),
    .A3(_01724_),
    .A4(_01732_),
    .ZN(_01733_));
 XNOR2_X1 _24925_ (.A(_01731_),
    .B(_01733_),
    .ZN(_01734_));
 INV_X1 _24926_ (.A(_21543_),
    .ZN(_01735_));
 INV_X1 _24927_ (.A(_21544_),
    .ZN(_01736_));
 OAI21_X1 _24928_ (.A(_01735_),
    .B1(_01736_),
    .B2(_14102_),
    .ZN(_01737_));
 AOI21_X1 _24929_ (.A(_21550_),
    .B1(_01737_),
    .B2(_21551_),
    .ZN(_01738_));
 XNOR2_X1 _24930_ (.A(_21555_),
    .B(_01738_),
    .ZN(_01739_));
 MUX2_X1 _24931_ (.A(_01734_),
    .B(_01739_),
    .S(_01597_),
    .Z(_01740_));
 NAND2_X1 _24932_ (.A1(_01418_),
    .A2(_21542_),
    .ZN(_01741_));
 OAI21_X1 _24933_ (.A(_01741_),
    .B1(_01732_),
    .B2(_01418_),
    .ZN(_01742_));
 MUX2_X1 _24934_ (.A(_14101_),
    .B(_01742_),
    .S(_01434_),
    .Z(_21545_));
 NAND3_X1 _24935_ (.A1(_21538_),
    .A2(_01728_),
    .A3(_21545_),
    .ZN(_01743_));
 XNOR2_X1 _24936_ (.A(_01740_),
    .B(_01743_),
    .ZN(_01744_));
 MUX2_X1 _24937_ (.A(\g_reduce0[2].adder.a[13] ),
    .B(_01744_),
    .S(_00956_),
    .Z(_01745_));
 MUX2_X2 _24938_ (.A(\g_reduce0[2].adder.b[13] ),
    .B(_01745_),
    .S(_01441_),
    .Z(_00068_));
 OR2_X1 _24939_ (.A1(_00953_),
    .A2(_01004_),
    .ZN(_01746_));
 NAND2_X1 _24940_ (.A1(\g_reduce0[2].adder.a[14] ),
    .A2(_01746_),
    .ZN(_01747_));
 NOR4_X1 _24941_ (.A1(_01597_),
    .A2(_01724_),
    .A3(_01725_),
    .A4(_01731_),
    .ZN(_01748_));
 AOI21_X1 _24942_ (.A(_21550_),
    .B1(_21551_),
    .B2(_14100_),
    .ZN(_01749_));
 INV_X1 _24943_ (.A(_01749_),
    .ZN(_01750_));
 AOI21_X1 _24944_ (.A(_21554_),
    .B1(_01750_),
    .B2(_21555_),
    .ZN(_01751_));
 AOI21_X1 _24945_ (.A(_01748_),
    .B1(_01751_),
    .B2(_01597_),
    .ZN(_01752_));
 NAND3_X1 _24946_ (.A1(_21546_),
    .A2(_01728_),
    .A3(_01740_),
    .ZN(_01753_));
 XNOR2_X2 _24947_ (.A(_01752_),
    .B(_01753_),
    .ZN(_01754_));
 MUX2_X1 _24948_ (.A(_01747_),
    .B(_01746_),
    .S(_01754_),
    .Z(_01755_));
 OAI22_X2 _24949_ (.A1(_00953_),
    .A2(_01441_),
    .B1(_01663_),
    .B2(_01755_),
    .ZN(_01756_));
 NOR2_X1 _24950_ (.A1(\g_reduce0[2].adder.a[14] ),
    .A2(_00951_),
    .ZN(_01757_));
 AOI21_X1 _24951_ (.A(_01663_),
    .B1(_01004_),
    .B2(_01754_),
    .ZN(_01758_));
 NAND2_X1 _24952_ (.A1(_00953_),
    .A2(_00973_),
    .ZN(_01759_));
 OAI21_X2 _24953_ (.A(_01758_),
    .B1(_01759_),
    .B2(_01754_),
    .ZN(_01760_));
 AOI21_X4 _24954_ (.A(_01756_),
    .B1(_01757_),
    .B2(_01760_),
    .ZN(_00069_));
 BUF_X2 _24955_ (.A(\g_reduce0[4].adder.a[12] ),
    .Z(_01761_));
 OR2_X1 _24956_ (.A1(\g_reduce0[4].adder.a[10] ),
    .A2(\g_reduce0[4].adder.a[13] ),
    .ZN(_01762_));
 OR4_X1 _24957_ (.A1(\g_reduce0[4].adder.a[11] ),
    .A2(_01761_),
    .A3(\g_reduce0[4].adder.a[14] ),
    .A4(_01762_),
    .ZN(_01763_));
 BUF_X4 _24958_ (.A(_01763_),
    .Z(_01764_));
 BUF_X2 _24959_ (.A(\g_reduce0[4].adder.b[12] ),
    .Z(_01765_));
 CLKBUF_X2 _24960_ (.A(\g_reduce0[4].adder.b[14] ),
    .Z(_01766_));
 OR2_X1 _24961_ (.A1(\g_reduce0[4].adder.b[10] ),
    .A2(\g_reduce0[4].adder.b[13] ),
    .ZN(_01767_));
 NOR4_X4 _24962_ (.A1(\g_reduce0[4].adder.b[11] ),
    .A2(_01765_),
    .A3(_01766_),
    .A4(_01767_),
    .ZN(_01768_));
 INV_X2 _24963_ (.A(_21599_),
    .ZN(_01769_));
 INV_X1 _24964_ (.A(_21560_),
    .ZN(_01770_));
 INV_X1 _24965_ (.A(_21566_),
    .ZN(_01771_));
 BUF_X2 _24966_ (.A(_21564_),
    .Z(_01772_));
 AOI21_X1 _24967_ (.A(_21563_),
    .B1(_01771_),
    .B2(_01772_),
    .ZN(_01773_));
 BUF_X4 _24968_ (.A(_21561_),
    .Z(_01774_));
 INV_X2 _24969_ (.A(_01774_),
    .ZN(_01775_));
 OAI21_X1 _24970_ (.A(_01770_),
    .B1(_01773_),
    .B2(_01775_),
    .ZN(_01776_));
 BUF_X2 _24971_ (.A(_21558_),
    .Z(_01777_));
 AOI21_X2 _24972_ (.A(_21557_),
    .B1(_01776_),
    .B2(_01777_),
    .ZN(_01778_));
 BUF_X2 _24973_ (.A(_21600_),
    .Z(_01779_));
 INV_X4 _24974_ (.A(_01779_),
    .ZN(_01780_));
 OAI21_X4 _24975_ (.A(_01769_),
    .B1(_01778_),
    .B2(_01780_),
    .ZN(_01781_));
 NAND4_X2 _24976_ (.A1(_21570_),
    .A2(_21573_),
    .A3(_21576_),
    .A4(_21579_),
    .ZN(_01782_));
 NAND3_X1 _24977_ (.A1(_21585_),
    .A2(_21588_),
    .A3(_21591_),
    .ZN(_01783_));
 INV_X1 _24978_ (.A(\g_reduce0[4].adder.a[0] ),
    .ZN(_01784_));
 OAI21_X1 _24979_ (.A(_21594_),
    .B1(\g_reduce0[4].adder.b[0] ),
    .B2(_01784_),
    .ZN(_01785_));
 INV_X1 _24980_ (.A(_21593_),
    .ZN(_01786_));
 AOI21_X1 _24981_ (.A(_01783_),
    .B1(_01785_),
    .B2(_01786_),
    .ZN(_01787_));
 INV_X1 _24982_ (.A(_21584_),
    .ZN(_01788_));
 AOI21_X1 _24983_ (.A(_21587_),
    .B1(_21588_),
    .B2(_21590_),
    .ZN(_01789_));
 INV_X1 _24984_ (.A(_21585_),
    .ZN(_01790_));
 OAI21_X1 _24985_ (.A(_01788_),
    .B1(_01789_),
    .B2(_01790_),
    .ZN(_01791_));
 OAI21_X2 _24986_ (.A(_21582_),
    .B1(_01787_),
    .B2(_01791_),
    .ZN(_01792_));
 INV_X1 _24987_ (.A(_21581_),
    .ZN(_01793_));
 AOI21_X4 _24988_ (.A(_01782_),
    .B1(_01792_),
    .B2(_01793_),
    .ZN(_01794_));
 INV_X1 _24989_ (.A(_21573_),
    .ZN(_01795_));
 AOI21_X1 _24990_ (.A(_21575_),
    .B1(_21576_),
    .B2(_21578_),
    .ZN(_01796_));
 NOR2_X1 _24991_ (.A1(_01795_),
    .A2(_01796_),
    .ZN(_01797_));
 OAI21_X2 _24992_ (.A(_21570_),
    .B1(_21572_),
    .B2(_01797_),
    .ZN(_01798_));
 CLKBUF_X3 _24993_ (.A(_21567_),
    .Z(_01799_));
 INV_X1 _24994_ (.A(_01799_),
    .ZN(_01800_));
 INV_X2 _24995_ (.A(_01777_),
    .ZN(_01801_));
 NOR4_X4 _24996_ (.A1(_01780_),
    .A2(_21569_),
    .A3(_01800_),
    .A4(_01801_),
    .ZN(_01802_));
 NAND4_X4 _24997_ (.A1(_01774_),
    .A2(_01772_),
    .A3(_01798_),
    .A4(_01802_),
    .ZN(_01803_));
 OAI21_X1 _24998_ (.A(_01781_),
    .B1(_01794_),
    .B2(_01803_),
    .ZN(_01804_));
 BUF_X1 _24999_ (.A(_01804_),
    .Z(_01805_));
 OAI21_X1 _25000_ (.A(_01764_),
    .B1(_01768_),
    .B2(_01805_),
    .ZN(_01806_));
 MUX2_X2 _25001_ (.A(\g_reduce0[4].adder.a[15] ),
    .B(\g_reduce0[4].adder.b[15] ),
    .S(_01806_),
    .Z(_00086_));
 OR2_X1 _25002_ (.A1(_01780_),
    .A2(_01778_),
    .ZN(_01807_));
 AND4_X1 _25003_ (.A1(_21570_),
    .A2(_21573_),
    .A3(_21576_),
    .A4(_21579_),
    .ZN(_01808_));
 INV_X1 _25004_ (.A(_21582_),
    .ZN(_01809_));
 AND3_X1 _25005_ (.A1(_21585_),
    .A2(_21588_),
    .A3(_21591_),
    .ZN(_01810_));
 INV_X1 _25006_ (.A(_21594_),
    .ZN(_01811_));
 INV_X1 _25007_ (.A(\g_reduce0[4].adder.b[0] ),
    .ZN(_01812_));
 AOI21_X1 _25008_ (.A(_01811_),
    .B1(_01812_),
    .B2(\g_reduce0[4].adder.a[0] ),
    .ZN(_01813_));
 OAI21_X1 _25009_ (.A(_01810_),
    .B1(_01813_),
    .B2(_21593_),
    .ZN(_01814_));
 INV_X1 _25010_ (.A(_01789_),
    .ZN(_01815_));
 AOI21_X1 _25011_ (.A(_21584_),
    .B1(_01815_),
    .B2(_21585_),
    .ZN(_01816_));
 AOI21_X1 _25012_ (.A(_01809_),
    .B1(_01814_),
    .B2(_01816_),
    .ZN(_01817_));
 OAI21_X2 _25013_ (.A(_01808_),
    .B1(_01817_),
    .B2(_21581_),
    .ZN(_01818_));
 AND4_X1 _25014_ (.A1(_01774_),
    .A2(_01772_),
    .A3(_01798_),
    .A4(_01802_),
    .ZN(_01819_));
 AOI22_X4 _25015_ (.A1(_01769_),
    .A2(_01807_),
    .B1(_01818_),
    .B2(_01819_),
    .ZN(_01820_));
 BUF_X4 _25016_ (.A(_01820_),
    .Z(_01821_));
 MUX2_X1 _25017_ (.A(\g_reduce0[4].adder.a[10] ),
    .B(\g_reduce0[4].adder.b[10] ),
    .S(_01821_),
    .Z(_21684_));
 NOR2_X1 _25018_ (.A1(\g_reduce0[4].adder.a[13] ),
    .A2(_00531_),
    .ZN(_01822_));
 NOR2_X1 _25019_ (.A1(\g_reduce0[4].adder.b[13] ),
    .A2(_21556_),
    .ZN(_01823_));
 MUX2_X1 _25020_ (.A(_01822_),
    .B(_01823_),
    .S(_01805_),
    .Z(_01824_));
 NOR2_X1 _25021_ (.A1(_01761_),
    .A2(_00528_),
    .ZN(_01825_));
 NOR2_X1 _25022_ (.A1(_01765_),
    .A2(_21559_),
    .ZN(_01826_));
 MUX2_X2 _25023_ (.A(_01825_),
    .B(_01826_),
    .S(_01804_),
    .Z(_01827_));
 NOR2_X1 _25024_ (.A1(\g_reduce0[4].adder.a[11] ),
    .A2(_00523_),
    .ZN(_01828_));
 OAI221_X2 _25025_ (.A(_01781_),
    .B1(_01794_),
    .B2(_01803_),
    .C1(_01828_),
    .C2(_21596_),
    .ZN(_01829_));
 NOR2_X2 _25026_ (.A1(\g_reduce0[4].adder.b[11] ),
    .A2(_21562_),
    .ZN(_01830_));
 NOR2_X2 _25027_ (.A1(_21596_),
    .A2(_01830_),
    .ZN(_01831_));
 OAI21_X2 _25028_ (.A(_01829_),
    .B1(_01831_),
    .B2(_01820_),
    .ZN(_01832_));
 OR4_X2 _25029_ (.A1(_01779_),
    .A2(_01824_),
    .A3(_01827_),
    .A4(_01832_),
    .ZN(_01833_));
 NOR2_X2 _25030_ (.A1(_01780_),
    .A2(_01801_),
    .ZN(_01834_));
 NOR3_X2 _25031_ (.A1(_01780_),
    .A2(_01801_),
    .A3(_01775_),
    .ZN(_01835_));
 AOI22_X4 _25032_ (.A1(_01827_),
    .A2(_01834_),
    .B1(_01835_),
    .B2(_01832_),
    .ZN(_01836_));
 OR4_X2 _25033_ (.A1(_01779_),
    .A2(_01774_),
    .A3(_01824_),
    .A4(_01827_),
    .ZN(_01837_));
 NAND2_X1 _25034_ (.A1(_01780_),
    .A2(_01801_),
    .ZN(_01838_));
 MUX2_X1 _25035_ (.A(_01838_),
    .B(_01780_),
    .S(_01824_),
    .Z(_01839_));
 NAND4_X4 _25036_ (.A1(_01833_),
    .A2(_01836_),
    .A3(_01837_),
    .A4(_01839_),
    .ZN(_01840_));
 OAI211_X2 _25037_ (.A(_01774_),
    .B(_01829_),
    .C1(_01831_),
    .C2(_01821_),
    .ZN(_01841_));
 NOR2_X1 _25038_ (.A1(_21596_),
    .A2(_01828_),
    .ZN(_01842_));
 OAI211_X4 _25039_ (.A(_01781_),
    .B(_01842_),
    .C1(_01803_),
    .C2(_01794_),
    .ZN(_01843_));
 OR2_X2 _25040_ (.A1(_21596_),
    .A2(_01830_),
    .ZN(_01844_));
 OAI211_X2 _25041_ (.A(_01775_),
    .B(_01843_),
    .C1(_01844_),
    .C2(_01820_),
    .ZN(_01845_));
 NAND2_X2 _25042_ (.A1(_01841_),
    .A2(_01845_),
    .ZN(_01846_));
 BUF_X4 _25043_ (.A(_01846_),
    .Z(_01847_));
 MUX2_X1 _25044_ (.A(_00518_),
    .B(_21592_),
    .S(_01821_),
    .Z(_01848_));
 CLKBUF_X3 _25045_ (.A(_01821_),
    .Z(_01849_));
 MUX2_X1 _25046_ (.A(_00519_),
    .B(_00520_),
    .S(_01849_),
    .Z(_01850_));
 CLKBUF_X3 _25047_ (.A(_01799_),
    .Z(_01851_));
 MUX2_X1 _25048_ (.A(_01848_),
    .B(_01850_),
    .S(_01851_),
    .Z(_01852_));
 MUX2_X1 _25049_ (.A(_00522_),
    .B(_21589_),
    .S(_01821_),
    .Z(_01853_));
 MUX2_X1 _25050_ (.A(_00521_),
    .B(_21586_),
    .S(_01849_),
    .Z(_01854_));
 CLKBUF_X3 _25051_ (.A(_01800_),
    .Z(_01855_));
 MUX2_X1 _25052_ (.A(_01853_),
    .B(_01854_),
    .S(_01855_),
    .Z(_01856_));
 BUF_X2 _25053_ (.A(_21597_),
    .Z(_01857_));
 CLKBUF_X3 _25054_ (.A(_01857_),
    .Z(_01858_));
 MUX2_X1 _25055_ (.A(_01852_),
    .B(_01856_),
    .S(_01858_),
    .Z(_01859_));
 BUF_X2 _25056_ (.A(_01858_),
    .Z(_01860_));
 NAND2_X1 _25057_ (.A1(_01855_),
    .A2(_01860_),
    .ZN(_01861_));
 MUX2_X1 _25058_ (.A(_00530_),
    .B(_21571_),
    .S(_01849_),
    .Z(_01862_));
 OR2_X1 _25059_ (.A1(_01855_),
    .A2(_01862_),
    .ZN(_01863_));
 MUX2_X1 _25060_ (.A(_00529_),
    .B(_21568_),
    .S(_01849_),
    .Z(_01864_));
 OAI21_X1 _25061_ (.A(_01863_),
    .B1(_01864_),
    .B2(_01851_),
    .ZN(_01865_));
 OAI21_X1 _25062_ (.A(_01861_),
    .B1(_01865_),
    .B2(_01860_),
    .ZN(_01866_));
 INV_X1 _25063_ (.A(\g_reduce0[4].adder.b[10] ),
    .ZN(_01867_));
 OR2_X1 _25064_ (.A1(\g_reduce0[4].adder.a[10] ),
    .A2(_01867_),
    .ZN(_01868_));
 AOI21_X1 _25065_ (.A(_01830_),
    .B1(_01868_),
    .B2(_01772_),
    .ZN(_01869_));
 OAI22_X1 _25066_ (.A1(_01765_),
    .A2(_21559_),
    .B1(_01775_),
    .B2(_01869_),
    .ZN(_01870_));
 AND2_X1 _25067_ (.A1(_01777_),
    .A2(_01870_),
    .ZN(_01871_));
 NOR2_X1 _25068_ (.A1(_01777_),
    .A2(_01870_),
    .ZN(_01872_));
 OAI21_X2 _25069_ (.A(_01805_),
    .B1(_01871_),
    .B2(_01872_),
    .ZN(_01873_));
 NAND2_X1 _25070_ (.A1(\g_reduce0[4].adder.a[10] ),
    .A2(_01867_),
    .ZN(_01874_));
 AOI21_X1 _25071_ (.A(_01828_),
    .B1(_01874_),
    .B2(_01772_),
    .ZN(_01875_));
 OAI22_X1 _25072_ (.A1(_01761_),
    .A2(_00528_),
    .B1(_01775_),
    .B2(_01875_),
    .ZN(_01876_));
 AND2_X1 _25073_ (.A1(_01777_),
    .A2(_01876_),
    .ZN(_01877_));
 NOR2_X1 _25074_ (.A1(_01777_),
    .A2(_01876_),
    .ZN(_01878_));
 OAI21_X2 _25075_ (.A(_01820_),
    .B1(_01877_),
    .B2(_01878_),
    .ZN(_01879_));
 AND2_X1 _25076_ (.A1(_01873_),
    .A2(_01879_),
    .ZN(_01880_));
 BUF_X4 _25077_ (.A(_01880_),
    .Z(_01881_));
 MUX2_X1 _25078_ (.A(_01859_),
    .B(_01866_),
    .S(_01881_),
    .Z(_01882_));
 NAND2_X4 _25079_ (.A1(_01873_),
    .A2(_01879_),
    .ZN(_01883_));
 NAND2_X1 _25080_ (.A1(_01883_),
    .A2(_01847_),
    .ZN(_01884_));
 MUX2_X1 _25081_ (.A(_00527_),
    .B(_21577_),
    .S(_01849_),
    .Z(_01885_));
 OR2_X1 _25082_ (.A1(_01855_),
    .A2(_01885_),
    .ZN(_01886_));
 MUX2_X1 _25083_ (.A(_00526_),
    .B(_21574_),
    .S(_01849_),
    .Z(_01887_));
 OAI21_X1 _25084_ (.A(_01886_),
    .B1(_01887_),
    .B2(_01851_),
    .ZN(_01888_));
 INV_X1 _25085_ (.A(_01888_),
    .ZN(_01889_));
 NAND2_X1 _25086_ (.A1(_01860_),
    .A2(_01889_),
    .ZN(_01890_));
 MUX2_X1 _25087_ (.A(_00525_),
    .B(_21583_),
    .S(_01821_),
    .Z(_01891_));
 OR2_X1 _25088_ (.A1(_01855_),
    .A2(_01891_),
    .ZN(_01892_));
 MUX2_X1 _25089_ (.A(_00524_),
    .B(_21580_),
    .S(_01849_),
    .Z(_01893_));
 OAI21_X1 _25090_ (.A(_01892_),
    .B1(_01893_),
    .B2(_01851_),
    .ZN(_01894_));
 OAI21_X1 _25091_ (.A(_01890_),
    .B1(_01894_),
    .B2(_01860_),
    .ZN(_01895_));
 OAI22_X1 _25092_ (.A1(_01847_),
    .A2(_01882_),
    .B1(_01884_),
    .B2(_01895_),
    .ZN(_01896_));
 NAND2_X1 _25093_ (.A1(_01840_),
    .A2(_01896_),
    .ZN(_21664_));
 INV_X1 _25094_ (.A(_21664_),
    .ZN(_21661_));
 AND4_X1 _25095_ (.A1(_01873_),
    .A2(_01879_),
    .A3(_01841_),
    .A4(_01845_),
    .ZN(_01897_));
 NAND2_X1 _25096_ (.A1(_01805_),
    .A2(_01823_),
    .ZN(_01898_));
 NOR2_X1 _25097_ (.A1(_01774_),
    .A2(_01826_),
    .ZN(_01899_));
 NOR2_X1 _25098_ (.A1(_01774_),
    .A2(_01825_),
    .ZN(_01900_));
 MUX2_X1 _25099_ (.A(_01899_),
    .B(_01900_),
    .S(_01820_),
    .Z(_01901_));
 OR2_X1 _25100_ (.A1(\g_reduce0[4].adder.a[13] ),
    .A2(_00531_),
    .ZN(_01902_));
 OAI221_X2 _25101_ (.A(_01898_),
    .B1(_01901_),
    .B2(_01801_),
    .C1(_01805_),
    .C2(_01902_),
    .ZN(_01903_));
 XNOR2_X2 _25102_ (.A(_01779_),
    .B(_01903_),
    .ZN(_01904_));
 BUF_X4 _25103_ (.A(_01904_),
    .Z(_01905_));
 AOI21_X1 _25104_ (.A(_01860_),
    .B1(_01864_),
    .B2(_01851_),
    .ZN(_01906_));
 AND3_X1 _25105_ (.A1(_01897_),
    .A2(_01905_),
    .A3(_01906_),
    .ZN(_01907_));
 NAND2_X1 _25106_ (.A1(_01840_),
    .A2(_01883_),
    .ZN(_01908_));
 NOR2_X1 _25107_ (.A1(_01855_),
    .A2(_01848_),
    .ZN(_01909_));
 NOR2_X1 _25108_ (.A1(_01851_),
    .A2(_01853_),
    .ZN(_01910_));
 NOR3_X1 _25109_ (.A1(_01858_),
    .A2(_01909_),
    .A3(_01910_),
    .ZN(_01911_));
 OAI211_X4 _25110_ (.A(_01775_),
    .B(_01829_),
    .C1(_01831_),
    .C2(_01820_),
    .ZN(_01912_));
 OAI211_X4 _25111_ (.A(_01774_),
    .B(_01843_),
    .C1(_01844_),
    .C2(_01820_),
    .ZN(_01913_));
 MUX2_X1 _25112_ (.A(_01891_),
    .B(_01854_),
    .S(_01851_),
    .Z(_01914_));
 AOI221_X2 _25113_ (.A(_01911_),
    .B1(_01912_),
    .B2(_01913_),
    .C1(_01858_),
    .C2(_01914_),
    .ZN(_01915_));
 NOR2_X1 _25114_ (.A1(_01855_),
    .A2(_01887_),
    .ZN(_01916_));
 NOR2_X1 _25115_ (.A1(_01851_),
    .A2(_01862_),
    .ZN(_01917_));
 OAI21_X1 _25116_ (.A(_01860_),
    .B1(_01916_),
    .B2(_01917_),
    .ZN(_01918_));
 MUX2_X1 _25117_ (.A(_01885_),
    .B(_01893_),
    .S(_01851_),
    .Z(_01919_));
 OAI21_X1 _25118_ (.A(_01918_),
    .B1(_01919_),
    .B2(_01860_),
    .ZN(_01920_));
 AOI21_X1 _25119_ (.A(_01915_),
    .B1(_01920_),
    .B2(_01847_),
    .ZN(_01921_));
 NOR2_X1 _25120_ (.A1(_01908_),
    .A2(_01921_),
    .ZN(_01922_));
 NOR2_X2 _25121_ (.A1(_01907_),
    .A2(_01922_),
    .ZN(_14109_));
 INV_X1 _25122_ (.A(_14109_),
    .ZN(_14104_));
 NOR2_X1 _25123_ (.A1(_01847_),
    .A2(_01908_),
    .ZN(_01923_));
 NAND2_X1 _25124_ (.A1(_01906_),
    .A2(_01923_),
    .ZN(_21616_));
 INV_X1 _25125_ (.A(_21616_),
    .ZN(_21620_));
 NAND2_X2 _25126_ (.A1(_01913_),
    .A2(_01912_),
    .ZN(_01924_));
 AND4_X2 _25127_ (.A1(_01833_),
    .A2(_01836_),
    .A3(_01837_),
    .A4(_01839_),
    .ZN(_01925_));
 NOR2_X1 _25128_ (.A1(_01925_),
    .A2(_01881_),
    .ZN(_01926_));
 NAND2_X1 _25129_ (.A1(_01924_),
    .A2(_01926_),
    .ZN(_01927_));
 OR2_X1 _25130_ (.A1(_01866_),
    .A2(_01927_),
    .ZN(_21609_));
 INV_X1 _25131_ (.A(_21609_),
    .ZN(_21613_));
 MUX2_X1 _25132_ (.A(_00526_),
    .B(_00529_),
    .S(_01858_),
    .Z(_01928_));
 NOR2_X1 _25133_ (.A1(_01799_),
    .A2(_01858_),
    .ZN(_01929_));
 AOI22_X1 _25134_ (.A1(_01851_),
    .A2(_01928_),
    .B1(_01929_),
    .B2(_00530_),
    .ZN(_01930_));
 MUX2_X1 _25135_ (.A(_21574_),
    .B(_21568_),
    .S(_01858_),
    .Z(_01931_));
 AOI22_X2 _25136_ (.A1(_21571_),
    .A2(_01929_),
    .B1(_01931_),
    .B2(_01799_),
    .ZN(_01932_));
 MUX2_X2 _25137_ (.A(_01930_),
    .B(_01932_),
    .S(_01821_),
    .Z(_01933_));
 NAND2_X1 _25138_ (.A1(_01923_),
    .A2(_01933_),
    .ZN(_21644_));
 INV_X1 _25139_ (.A(_21644_),
    .ZN(_21648_));
 MUX2_X1 _25140_ (.A(_01888_),
    .B(_01865_),
    .S(_01860_),
    .Z(_01934_));
 NOR2_X2 _25141_ (.A1(_01855_),
    .A2(_01858_),
    .ZN(_01935_));
 MUX2_X1 _25142_ (.A(_01934_),
    .B(_01935_),
    .S(_01847_),
    .Z(_01936_));
 NAND2_X1 _25143_ (.A1(_01926_),
    .A2(_01936_),
    .ZN(_21623_));
 INV_X1 _25144_ (.A(_21623_),
    .ZN(_21627_));
 MUX2_X1 _25145_ (.A(_01906_),
    .B(_01920_),
    .S(_01924_),
    .Z(_01937_));
 AND2_X1 _25146_ (.A1(_01926_),
    .A2(_01937_),
    .ZN(_21630_));
 INV_X1 _25147_ (.A(_21630_),
    .ZN(_21634_));
 MUX2_X1 _25148_ (.A(_01895_),
    .B(_01866_),
    .S(_01847_),
    .Z(_01938_));
 NOR2_X1 _25149_ (.A1(_01908_),
    .A2(_01938_),
    .ZN(_21637_));
 INV_X1 _25150_ (.A(_21637_),
    .ZN(_21641_));
 AND2_X1 _25151_ (.A1(_01805_),
    .A2(_01930_),
    .ZN(_01939_));
 AOI21_X1 _25152_ (.A(_01939_),
    .B1(_01932_),
    .B2(_01849_),
    .ZN(_01940_));
 MUX2_X1 _25153_ (.A(_21583_),
    .B(_21577_),
    .S(_01857_),
    .Z(_01941_));
 MUX2_X1 _25154_ (.A(_21586_),
    .B(_21580_),
    .S(_01857_),
    .Z(_01942_));
 MUX2_X1 _25155_ (.A(_01941_),
    .B(_01942_),
    .S(_01799_),
    .Z(_01943_));
 MUX2_X1 _25156_ (.A(_00525_),
    .B(_00527_),
    .S(_01857_),
    .Z(_01944_));
 MUX2_X1 _25157_ (.A(_00521_),
    .B(_00524_),
    .S(_01858_),
    .Z(_01945_));
 MUX2_X1 _25158_ (.A(_01944_),
    .B(_01945_),
    .S(_01799_),
    .Z(_01946_));
 MUX2_X2 _25159_ (.A(_01943_),
    .B(_01946_),
    .S(_01805_),
    .Z(_01947_));
 MUX2_X1 _25160_ (.A(_01940_),
    .B(_01947_),
    .S(_01924_),
    .Z(_01948_));
 NOR2_X1 _25161_ (.A1(_01908_),
    .A2(_01948_),
    .ZN(_21655_));
 INV_X1 _25162_ (.A(_21655_),
    .ZN(_21658_));
 NOR2_X1 _25163_ (.A1(_01881_),
    .A2(_01924_),
    .ZN(_01949_));
 NAND3_X1 _25164_ (.A1(_01860_),
    .A2(_01883_),
    .A3(_01894_),
    .ZN(_01950_));
 MUX2_X1 _25165_ (.A(_01855_),
    .B(_01856_),
    .S(_01883_),
    .Z(_01951_));
 OAI21_X1 _25166_ (.A(_01950_),
    .B1(_01951_),
    .B2(_01860_),
    .ZN(_01952_));
 AOI22_X1 _25167_ (.A1(_01949_),
    .A2(_01934_),
    .B1(_01952_),
    .B2(_01924_),
    .ZN(_01953_));
 OR2_X1 _25168_ (.A1(_01925_),
    .A2(_01953_),
    .ZN(_21651_));
 INV_X1 _25169_ (.A(_21651_),
    .ZN(_21605_));
 XOR2_X2 _25170_ (.A(\g_reduce0[4].adder.a[15] ),
    .B(\g_reduce0[4].adder.b[15] ),
    .Z(_01954_));
 BUF_X4 _25171_ (.A(_01954_),
    .Z(_01955_));
 BUF_X2 _25172_ (.A(_21612_),
    .Z(_01956_));
 INV_X1 _25173_ (.A(_01956_),
    .ZN(_01957_));
 BUF_X2 _25174_ (.A(_21647_),
    .Z(_01958_));
 INV_X1 _25175_ (.A(_01958_),
    .ZN(_01959_));
 INV_X1 _25176_ (.A(_21628_),
    .ZN(_01960_));
 CLKBUF_X2 _25177_ (.A(_21633_),
    .Z(_01961_));
 NOR2_X1 _25178_ (.A1(_01961_),
    .A2(_21632_),
    .ZN(_01962_));
 BUF_X2 _25179_ (.A(_21626_),
    .Z(_01963_));
 OAI21_X1 _25180_ (.A(_01960_),
    .B1(_01962_),
    .B2(_01963_),
    .ZN(_01964_));
 NOR3_X1 _25181_ (.A1(_21628_),
    .A2(_21632_),
    .A3(_21639_),
    .ZN(_01965_));
 INV_X1 _25182_ (.A(_21607_),
    .ZN(_01966_));
 INV_X1 _25183_ (.A(_21608_),
    .ZN(_01967_));
 AOI21_X1 _25184_ (.A(_21601_),
    .B1(_14103_),
    .B2(_21602_),
    .ZN(_01968_));
 OAI21_X1 _25185_ (.A(_01966_),
    .B1(_01967_),
    .B2(_01968_),
    .ZN(_01969_));
 CLKBUF_X2 _25186_ (.A(_21657_),
    .Z(_01970_));
 AOI21_X1 _25187_ (.A(_21656_),
    .B1(_01969_),
    .B2(_01970_),
    .ZN(_01971_));
 BUF_X2 _25188_ (.A(_21640_),
    .Z(_01972_));
 INV_X1 _25189_ (.A(_01972_),
    .ZN(_01973_));
 OAI21_X1 _25190_ (.A(_01965_),
    .B1(_01971_),
    .B2(_01973_),
    .ZN(_01974_));
 AND3_X1 _25191_ (.A1(_01959_),
    .A2(_01964_),
    .A3(_01974_),
    .ZN(_01975_));
 OAI21_X1 _25192_ (.A(_01957_),
    .B1(_01975_),
    .B2(_21649_),
    .ZN(_01976_));
 NOR2_X1 _25193_ (.A1(_21621_),
    .A2(_21614_),
    .ZN(_01977_));
 INV_X1 _25194_ (.A(_21621_),
    .ZN(_01978_));
 BUF_X2 _25195_ (.A(_21619_),
    .Z(_01979_));
 AOI221_X2 _25196_ (.A(_01955_),
    .B1(_01976_),
    .B2(_01977_),
    .C1(_01978_),
    .C2(_01979_),
    .ZN(_01980_));
 OR2_X2 _25197_ (.A1(_01855_),
    .A2(_01858_),
    .ZN(_01981_));
 XNOR2_X2 _25198_ (.A(\g_reduce0[4].adder.a[15] ),
    .B(\g_reduce0[4].adder.b[15] ),
    .ZN(_01982_));
 CLKBUF_X3 _25199_ (.A(_01982_),
    .Z(_01983_));
 BUF_X4 _25200_ (.A(_01983_),
    .Z(_01984_));
 INV_X1 _25201_ (.A(_21625_),
    .ZN(_01985_));
 INV_X1 _25202_ (.A(_21642_),
    .ZN(_01986_));
 AOI21_X2 _25203_ (.A(_01961_),
    .B1(_01972_),
    .B2(_01986_),
    .ZN(_01987_));
 OAI21_X2 _25204_ (.A(_01963_),
    .B1(_21635_),
    .B2(_01987_),
    .ZN(_01988_));
 NOR4_X2 _25205_ (.A1(_21635_),
    .A2(_21625_),
    .A3(_21642_),
    .A4(_21659_),
    .ZN(_01989_));
 INV_X2 _25206_ (.A(_01970_),
    .ZN(_01990_));
 INV_X1 _25207_ (.A(_21652_),
    .ZN(_01991_));
 INV_X1 _25208_ (.A(_21653_),
    .ZN(_01992_));
 AOI21_X1 _25209_ (.A(_21603_),
    .B1(_14108_),
    .B2(_21604_),
    .ZN(_01993_));
 OAI21_X2 _25210_ (.A(_01991_),
    .B1(_01992_),
    .B2(_01993_),
    .ZN(_01994_));
 NAND2_X1 _25211_ (.A1(_01990_),
    .A2(_01994_),
    .ZN(_01995_));
 AOI22_X4 _25212_ (.A1(_01985_),
    .A2(_01988_),
    .B1(_01989_),
    .B2(_01995_),
    .ZN(_01996_));
 AOI21_X1 _25213_ (.A(_21646_),
    .B1(_01996_),
    .B2(_01958_),
    .ZN(_01997_));
 NOR2_X1 _25214_ (.A1(_01957_),
    .A2(_01997_),
    .ZN(_01998_));
 OAI21_X2 _25215_ (.A(_01979_),
    .B1(_21611_),
    .B2(_01998_),
    .ZN(_01999_));
 INV_X1 _25216_ (.A(_21618_),
    .ZN(_02000_));
 AOI21_X4 _25217_ (.A(_01984_),
    .B1(_01999_),
    .B2(_02000_),
    .ZN(_02001_));
 NOR4_X4 _25218_ (.A1(_01881_),
    .A2(_01847_),
    .A3(_01981_),
    .A4(_02001_),
    .ZN(_02002_));
 AOI21_X4 _25219_ (.A(_01980_),
    .B1(_02002_),
    .B2(_01905_),
    .ZN(_02003_));
 OR3_X1 _25220_ (.A1(_21618_),
    .A2(_21611_),
    .A3(_01983_),
    .ZN(_02004_));
 AOI21_X1 _25221_ (.A(_21646_),
    .B1(_21625_),
    .B2(_01958_),
    .ZN(_02005_));
 NAND2_X1 _25222_ (.A1(_01963_),
    .A2(_01958_),
    .ZN(_02006_));
 NOR2_X1 _25223_ (.A1(_21642_),
    .A2(_21659_),
    .ZN(_02007_));
 AOI21_X2 _25224_ (.A(_21652_),
    .B1(_14110_),
    .B2(_21653_),
    .ZN(_02008_));
 OAI21_X1 _25225_ (.A(_02007_),
    .B1(_02008_),
    .B2(_01970_),
    .ZN(_02009_));
 AOI21_X1 _25226_ (.A(_21635_),
    .B1(_01987_),
    .B2(_02009_),
    .ZN(_02010_));
 OAI21_X1 _25227_ (.A(_02005_),
    .B1(_02006_),
    .B2(_02010_),
    .ZN(_02011_));
 AOI21_X1 _25228_ (.A(_02004_),
    .B1(_02011_),
    .B2(_01956_),
    .ZN(_02012_));
 AOI21_X1 _25229_ (.A(_01979_),
    .B1(_21618_),
    .B2(_01955_),
    .ZN(_02013_));
 NOR2_X1 _25230_ (.A1(_21614_),
    .A2(_01954_),
    .ZN(_02014_));
 AOI21_X1 _25231_ (.A(_01958_),
    .B1(_01960_),
    .B2(_01963_),
    .ZN(_02015_));
 NOR2_X1 _25232_ (.A1(_21628_),
    .A2(_21632_),
    .ZN(_02016_));
 INV_X1 _25233_ (.A(_21656_),
    .ZN(_02017_));
 AOI21_X1 _25234_ (.A(_21607_),
    .B1(_14106_),
    .B2(_21608_),
    .ZN(_02018_));
 OAI21_X1 _25235_ (.A(_02017_),
    .B1(_02018_),
    .B2(_01990_),
    .ZN(_02019_));
 AOI21_X1 _25236_ (.A(_21639_),
    .B1(_02019_),
    .B2(_01972_),
    .ZN(_02020_));
 INV_X1 _25237_ (.A(_01961_),
    .ZN(_02021_));
 OAI21_X1 _25238_ (.A(_02016_),
    .B1(_02020_),
    .B2(_02021_),
    .ZN(_02022_));
 AOI21_X1 _25239_ (.A(_21649_),
    .B1(_02015_),
    .B2(_02022_),
    .ZN(_02023_));
 OAI21_X1 _25240_ (.A(_02014_),
    .B1(_02023_),
    .B2(_01956_),
    .ZN(_02024_));
 AOI221_X1 _25241_ (.A(_02012_),
    .B1(_02013_),
    .B2(_02024_),
    .C1(_21621_),
    .C2(_01984_),
    .ZN(_02025_));
 NAND3_X4 _25242_ (.A1(_01883_),
    .A2(_01924_),
    .A3(_01935_),
    .ZN(_02026_));
 XNOR2_X2 _25243_ (.A(_01780_),
    .B(_01903_),
    .ZN(_02027_));
 OAI21_X4 _25244_ (.A(_02025_),
    .B1(_02026_),
    .B2(_02027_),
    .ZN(_02028_));
 NOR3_X4 _25245_ (.A1(_01881_),
    .A2(_01846_),
    .A3(_01981_),
    .ZN(_02029_));
 INV_X2 _25246_ (.A(_02025_),
    .ZN(_02030_));
 NAND3_X4 _25247_ (.A1(_01904_),
    .A2(_02029_),
    .A3(_02030_),
    .ZN(_02031_));
 INV_X1 _25248_ (.A(_21649_),
    .ZN(_02032_));
 OAI21_X2 _25249_ (.A(_02014_),
    .B1(_01956_),
    .B2(_02032_),
    .ZN(_02033_));
 OR3_X1 _25250_ (.A1(_21646_),
    .A2(_21611_),
    .A3(_01982_),
    .ZN(_02034_));
 AOI21_X2 _25251_ (.A(_02034_),
    .B1(_01996_),
    .B2(_01958_),
    .ZN(_02035_));
 OAI21_X1 _25252_ (.A(_01983_),
    .B1(_21614_),
    .B2(_01957_),
    .ZN(_02036_));
 OAI21_X2 _25253_ (.A(_02036_),
    .B1(_21611_),
    .B2(_01956_),
    .ZN(_02037_));
 OAI22_X4 _25254_ (.A1(_01975_),
    .A2(_02033_),
    .B1(_02035_),
    .B2(_02037_),
    .ZN(_02038_));
 XOR2_X2 _25255_ (.A(_01979_),
    .B(_02038_),
    .Z(_02039_));
 MUX2_X2 _25256_ (.A(_02023_),
    .B(_02011_),
    .S(_01955_),
    .Z(_02040_));
 XNOR2_X2 _25257_ (.A(_01956_),
    .B(_02040_),
    .ZN(_02041_));
 NOR2_X1 _25258_ (.A1(_01958_),
    .A2(_01983_),
    .ZN(_02042_));
 NOR2_X1 _25259_ (.A1(_01959_),
    .A2(_01983_),
    .ZN(_02043_));
 MUX2_X1 _25260_ (.A(_02042_),
    .B(_02043_),
    .S(_01996_),
    .Z(_02044_));
 AND4_X1 _25261_ (.A1(_01959_),
    .A2(_01964_),
    .A3(_01974_),
    .A4(_01984_),
    .ZN(_02045_));
 NAND2_X1 _25262_ (.A1(_01958_),
    .A2(_01984_),
    .ZN(_02046_));
 AOI21_X2 _25263_ (.A(_02046_),
    .B1(_01974_),
    .B2(_01964_),
    .ZN(_02047_));
 OR3_X2 _25264_ (.A1(_02044_),
    .A2(_02045_),
    .A3(_02047_),
    .ZN(_02048_));
 INV_X1 _25265_ (.A(_21632_),
    .ZN(_02049_));
 OAI21_X1 _25266_ (.A(_02049_),
    .B1(_02020_),
    .B2(_02021_),
    .ZN(_02050_));
 MUX2_X2 _25267_ (.A(_02010_),
    .B(_02050_),
    .S(_01983_),
    .Z(_02051_));
 XNOR2_X2 _25268_ (.A(_01963_),
    .B(_02051_),
    .ZN(_02052_));
 AOI21_X1 _25269_ (.A(_01982_),
    .B1(_01986_),
    .B2(_01972_),
    .ZN(_02053_));
 AOI21_X1 _25270_ (.A(_21639_),
    .B1(_21656_),
    .B2(_01972_),
    .ZN(_02054_));
 AOI21_X2 _25271_ (.A(_02053_),
    .B1(_01983_),
    .B2(_02054_),
    .ZN(_02055_));
 NAND2_X1 _25272_ (.A1(_01954_),
    .A2(_02007_),
    .ZN(_02056_));
 AOI21_X2 _25273_ (.A(_02056_),
    .B1(_01994_),
    .B2(_01990_),
    .ZN(_02057_));
 AND4_X1 _25274_ (.A1(_01972_),
    .A2(_01970_),
    .A3(_01969_),
    .A4(_01982_),
    .ZN(_02058_));
 NOR3_X4 _25275_ (.A1(_02055_),
    .A2(_02057_),
    .A3(_02058_),
    .ZN(_02059_));
 XNOR2_X2 _25276_ (.A(_01961_),
    .B(_02059_),
    .ZN(_02060_));
 NOR2_X1 _25277_ (.A1(_01954_),
    .A2(_02019_),
    .ZN(_02061_));
 INV_X1 _25278_ (.A(_21659_),
    .ZN(_02062_));
 OAI21_X2 _25279_ (.A(_02062_),
    .B1(_02008_),
    .B2(_01970_),
    .ZN(_02063_));
 AOI21_X4 _25280_ (.A(_02061_),
    .B1(_02063_),
    .B2(_01955_),
    .ZN(_02064_));
 XNOR2_X2 _25281_ (.A(_01972_),
    .B(_02064_),
    .ZN(_02065_));
 AND2_X1 _25282_ (.A1(_01969_),
    .A2(_01983_),
    .ZN(_02066_));
 NOR2_X1 _25283_ (.A1(_01983_),
    .A2(_01994_),
    .ZN(_02067_));
 OR3_X2 _25284_ (.A1(_01990_),
    .A2(_02066_),
    .A3(_02067_),
    .ZN(_02068_));
 OAI21_X2 _25285_ (.A(_01990_),
    .B1(_02066_),
    .B2(_02067_),
    .ZN(_02069_));
 XOR2_X1 _25286_ (.A(_14106_),
    .B(_21608_),
    .Z(_02070_));
 NAND2_X1 _25287_ (.A1(_01982_),
    .A2(_02070_),
    .ZN(_02071_));
 XOR2_X1 _25288_ (.A(_14110_),
    .B(_21653_),
    .Z(_02072_));
 NAND2_X1 _25289_ (.A1(_01954_),
    .A2(_02072_),
    .ZN(_02073_));
 AND2_X1 _25290_ (.A1(_02071_),
    .A2(_02073_),
    .ZN(_02074_));
 BUF_X2 _25291_ (.A(_02074_),
    .Z(_02075_));
 INV_X1 _25292_ (.A(_14111_),
    .ZN(_02076_));
 INV_X1 _25293_ (.A(_14107_),
    .ZN(_02077_));
 MUX2_X2 _25294_ (.A(_02076_),
    .B(_02077_),
    .S(_01983_),
    .Z(_02078_));
 NAND2_X1 _25295_ (.A1(_02075_),
    .A2(_02078_),
    .ZN(_02079_));
 NAND3_X1 _25296_ (.A1(_02068_),
    .A2(_02069_),
    .A3(_02079_),
    .ZN(_02080_));
 AOI21_X1 _25297_ (.A(_02060_),
    .B1(_02065_),
    .B2(_02080_),
    .ZN(_02081_));
 OAI21_X2 _25298_ (.A(_02048_),
    .B1(_02052_),
    .B2(_02081_),
    .ZN(_02082_));
 AOI21_X4 _25299_ (.A(_02039_),
    .B1(_02041_),
    .B2(_02082_),
    .ZN(_02083_));
 XOR2_X2 _25300_ (.A(_01963_),
    .B(_02051_),
    .Z(_02084_));
 NAND2_X4 _25301_ (.A1(_02071_),
    .A2(_02073_),
    .ZN(_02085_));
 MUX2_X1 _25302_ (.A(_21663_),
    .B(_21665_),
    .S(_01955_),
    .Z(_02086_));
 NOR2_X1 _25303_ (.A1(_02085_),
    .A2(_02086_),
    .ZN(_02087_));
 NAND4_X2 _25304_ (.A1(_02041_),
    .A2(_02084_),
    .A3(_02065_),
    .A4(_02087_),
    .ZN(_02088_));
 NAND2_X2 _25305_ (.A1(_02083_),
    .A2(_02088_),
    .ZN(_02089_));
 NAND3_X4 _25306_ (.A1(_02028_),
    .A2(_02031_),
    .A3(_02089_),
    .ZN(_02090_));
 XNOR2_X2 _25307_ (.A(_01979_),
    .B(_02038_),
    .ZN(_02091_));
 XNOR2_X2 _25308_ (.A(_01957_),
    .B(_02040_),
    .ZN(_02092_));
 NOR3_X2 _25309_ (.A1(_02044_),
    .A2(_02045_),
    .A3(_02047_),
    .ZN(_02093_));
 XNOR2_X2 _25310_ (.A(_02021_),
    .B(_02059_),
    .ZN(_02094_));
 XNOR2_X2 _25311_ (.A(_01973_),
    .B(_02064_),
    .ZN(_02095_));
 AND3_X1 _25312_ (.A1(_02068_),
    .A2(_02069_),
    .A3(_02079_),
    .ZN(_02096_));
 OAI21_X1 _25313_ (.A(_02094_),
    .B1(_02095_),
    .B2(_02096_),
    .ZN(_02097_));
 AOI21_X2 _25314_ (.A(_02093_),
    .B1(_02084_),
    .B2(_02097_),
    .ZN(_02098_));
 OAI21_X4 _25315_ (.A(_02091_),
    .B1(_02092_),
    .B2(_02098_),
    .ZN(_02099_));
 NAND3_X2 _25316_ (.A1(_01913_),
    .A2(_01912_),
    .A3(_01947_),
    .ZN(_02100_));
 MUX2_X1 _25317_ (.A(_00519_),
    .B(_00522_),
    .S(_01857_),
    .Z(_02101_));
 NOR2_X1 _25318_ (.A1(_01799_),
    .A2(_02101_),
    .ZN(_02102_));
 MUX2_X1 _25319_ (.A(_00520_),
    .B(_21589_),
    .S(_01857_),
    .Z(_02103_));
 NOR2_X1 _25320_ (.A1(_01799_),
    .A2(_02103_),
    .ZN(_02104_));
 MUX2_X1 _25321_ (.A(_02102_),
    .B(_02104_),
    .S(_01820_),
    .Z(_02105_));
 NAND2_X1 _25322_ (.A1(_01799_),
    .A2(_01857_),
    .ZN(_02106_));
 NOR2_X1 _25323_ (.A1(_00518_),
    .A2(_02106_),
    .ZN(_02107_));
 NOR2_X1 _25324_ (.A1(_21592_),
    .A2(_02106_),
    .ZN(_02108_));
 MUX2_X1 _25325_ (.A(_02107_),
    .B(_02108_),
    .S(_01820_),
    .Z(_02109_));
 OR2_X1 _25326_ (.A1(_02105_),
    .A2(_02109_),
    .ZN(_02110_));
 OAI211_X4 _25327_ (.A(_01883_),
    .B(_02100_),
    .C1(_02110_),
    .C2(_01847_),
    .ZN(_02111_));
 AOI21_X2 _25328_ (.A(_01955_),
    .B1(_01933_),
    .B2(_01897_),
    .ZN(_02112_));
 AOI22_X4 _25329_ (.A1(_01925_),
    .A2(_01984_),
    .B1(_02111_),
    .B2(_02112_),
    .ZN(_02113_));
 NAND3_X1 _25330_ (.A1(_01873_),
    .A2(_01879_),
    .A3(_01933_),
    .ZN(_02114_));
 NOR2_X1 _25331_ (.A1(_01847_),
    .A2(_02114_),
    .ZN(_02115_));
 AOI211_X2 _25332_ (.A(_02105_),
    .B(_02109_),
    .C1(_01913_),
    .C2(_01912_),
    .ZN(_02116_));
 AOI211_X2 _25333_ (.A(_01881_),
    .B(_02116_),
    .C1(_01947_),
    .C2(_01846_),
    .ZN(_02117_));
 OAI211_X2 _25334_ (.A(_01840_),
    .B(_01955_),
    .C1(_02115_),
    .C2(_02117_),
    .ZN(_02118_));
 AOI21_X4 _25335_ (.A(_02099_),
    .B1(_02113_),
    .B2(_02118_),
    .ZN(_02119_));
 OAI21_X4 _25336_ (.A(_02003_),
    .B1(_02090_),
    .B2(_02119_),
    .ZN(_21666_));
 INV_X4 _25337_ (.A(_21666_),
    .ZN(_21669_));
 INV_X1 _25338_ (.A(_21672_),
    .ZN(_02120_));
 INV_X1 _25339_ (.A(_01980_),
    .ZN(_02121_));
 NAND2_X1 _25340_ (.A1(_02121_),
    .A2(_02030_),
    .ZN(_02122_));
 NAND2_X2 _25341_ (.A1(_02048_),
    .A2(_02084_),
    .ZN(_02123_));
 NOR3_X4 _25342_ (.A1(_02039_),
    .A2(_02092_),
    .A3(_02123_),
    .ZN(_02124_));
 AND2_X2 _25343_ (.A1(_02068_),
    .A2(_02069_),
    .ZN(_02125_));
 NAND2_X1 _25344_ (.A1(_02125_),
    .A2(_02075_),
    .ZN(_02126_));
 NAND2_X1 _25345_ (.A1(_02094_),
    .A2(_02065_),
    .ZN(_02127_));
 OR2_X2 _25346_ (.A1(_02126_),
    .A2(_02127_),
    .ZN(_02128_));
 AOI221_X2 _25347_ (.A(_02122_),
    .B1(_02124_),
    .B2(_02128_),
    .C1(_01905_),
    .C2(_02029_),
    .ZN(_02129_));
 NAND2_X1 _25348_ (.A1(_02128_),
    .A2(_02124_),
    .ZN(_02130_));
 AND2_X1 _25349_ (.A1(_02001_),
    .A2(_02025_),
    .ZN(_02131_));
 AND4_X2 _25350_ (.A1(_01905_),
    .A2(_02029_),
    .A3(_02130_),
    .A4(_02131_),
    .ZN(_02132_));
 NOR3_X4 _25351_ (.A1(_02120_),
    .A2(_02129_),
    .A3(_02132_),
    .ZN(_02133_));
 NOR2_X2 _25352_ (.A1(_01980_),
    .A2(_02025_),
    .ZN(_02134_));
 INV_X1 _25353_ (.A(_02124_),
    .ZN(_02135_));
 INV_X1 _25354_ (.A(_02128_),
    .ZN(_02136_));
 OAI221_X2 _25355_ (.A(_02134_),
    .B1(_02135_),
    .B2(_02136_),
    .C1(_02027_),
    .C2(_02026_),
    .ZN(_02137_));
 NAND4_X4 _25356_ (.A1(_01905_),
    .A2(_02029_),
    .A3(_02130_),
    .A4(_02131_),
    .ZN(_02138_));
 AOI21_X4 _25357_ (.A(_21672_),
    .B1(_02137_),
    .B2(_02138_),
    .ZN(_02139_));
 NOR2_X2 _25358_ (.A1(_02133_),
    .A2(_02139_),
    .ZN(_02140_));
 INV_X1 _25359_ (.A(_02140_),
    .ZN(_02141_));
 CLKBUF_X3 _25360_ (.A(_02141_),
    .Z(_21692_));
 AOI21_X2 _25361_ (.A(_02122_),
    .B1(_02029_),
    .B2(_01905_),
    .ZN(_02142_));
 AND3_X1 _25362_ (.A1(_01905_),
    .A2(_02029_),
    .A3(_02131_),
    .ZN(_02143_));
 NOR2_X2 _25363_ (.A1(_02142_),
    .A2(_02143_),
    .ZN(_02144_));
 BUF_X4 _25364_ (.A(_02144_),
    .Z(_02145_));
 OAI21_X1 _25365_ (.A(_02124_),
    .B1(_02142_),
    .B2(_02143_),
    .ZN(_02146_));
 NOR3_X1 _25366_ (.A1(_02077_),
    .A2(_21663_),
    .A3(_01955_),
    .ZN(_02147_));
 NOR3_X1 _25367_ (.A1(_02076_),
    .A2(_21665_),
    .A3(_01984_),
    .ZN(_02148_));
 NOR3_X1 _25368_ (.A1(_02126_),
    .A2(_02147_),
    .A3(_02148_),
    .ZN(_02149_));
 NOR2_X1 _25369_ (.A1(_02127_),
    .A2(_02149_),
    .ZN(_02150_));
 AND2_X1 _25370_ (.A1(_02083_),
    .A2(_02150_),
    .ZN(_02151_));
 OAI211_X2 _25371_ (.A(_02124_),
    .B(_02151_),
    .C1(_02143_),
    .C2(_02142_),
    .ZN(_02152_));
 OAI21_X2 _25372_ (.A(_01984_),
    .B1(_02114_),
    .B2(_01847_),
    .ZN(_02153_));
 OAI22_X4 _25373_ (.A1(_01840_),
    .A2(_01955_),
    .B1(_02117_),
    .B2(_02153_),
    .ZN(_02154_));
 NAND2_X1 _25374_ (.A1(_01897_),
    .A2(_01933_),
    .ZN(_02155_));
 AOI211_X2 _25375_ (.A(_01925_),
    .B(_01984_),
    .C1(_02155_),
    .C2(_02111_),
    .ZN(_02156_));
 NOR3_X1 _25376_ (.A1(_02154_),
    .A2(_02156_),
    .A3(_02088_),
    .ZN(_02157_));
 OAI221_X2 _25377_ (.A(_02003_),
    .B1(_02128_),
    .B2(_02146_),
    .C1(_02152_),
    .C2(_02157_),
    .ZN(_02158_));
 BUF_X4 _25378_ (.A(_02158_),
    .Z(_02159_));
 NOR2_X2 _25379_ (.A1(_02145_),
    .A2(_02159_),
    .ZN(_02160_));
 BUF_X1 _25380_ (.A(_14112_),
    .Z(_02161_));
 INV_X1 _25381_ (.A(_02161_),
    .ZN(_02162_));
 BUF_X4 _25382_ (.A(_02162_),
    .Z(_02163_));
 OAI21_X4 _25383_ (.A(_02003_),
    .B1(_02133_),
    .B2(_02139_),
    .ZN(_02164_));
 NOR2_X4 _25384_ (.A1(_02154_),
    .A2(_02156_),
    .ZN(_02165_));
 NOR2_X1 _25385_ (.A1(_02025_),
    .A2(_02083_),
    .ZN(_02166_));
 OAI21_X1 _25386_ (.A(_02166_),
    .B1(_02026_),
    .B2(_02027_),
    .ZN(_02167_));
 NAND4_X2 _25387_ (.A1(_01905_),
    .A2(_02029_),
    .A3(_02025_),
    .A4(_02099_),
    .ZN(_02168_));
 NAND2_X2 _25388_ (.A1(_02167_),
    .A2(_02168_),
    .ZN(_02169_));
 NOR2_X2 _25389_ (.A1(_02165_),
    .A2(_02169_),
    .ZN(_02170_));
 NOR3_X4 _25390_ (.A1(_02163_),
    .A2(_02164_),
    .A3(_02170_),
    .ZN(_02171_));
 BUF_X2 _25391_ (.A(_21668_),
    .Z(_02172_));
 INV_X2 _25392_ (.A(_02172_),
    .ZN(_02173_));
 BUF_X4 _25393_ (.A(_02173_),
    .Z(_02174_));
 OAI21_X2 _25394_ (.A(_02174_),
    .B1(_02154_),
    .B2(_02156_),
    .ZN(_02175_));
 AOI22_X4 _25395_ (.A1(_02160_),
    .A2(_02171_),
    .B1(_02175_),
    .B2(_02145_),
    .ZN(_02176_));
 OAI21_X2 _25396_ (.A(_02134_),
    .B1(_02026_),
    .B2(_02027_),
    .ZN(_02177_));
 NAND3_X2 _25397_ (.A1(_01905_),
    .A2(_02029_),
    .A3(_02131_),
    .ZN(_02178_));
 NAND2_X4 _25398_ (.A1(_02177_),
    .A2(_02178_),
    .ZN(_02179_));
 BUF_X4 _25399_ (.A(_02179_),
    .Z(_02180_));
 NOR2_X1 _25400_ (.A1(_02174_),
    .A2(_02180_),
    .ZN(_02181_));
 AND2_X1 _25401_ (.A1(_21663_),
    .A2(_01984_),
    .ZN(_02182_));
 AOI21_X4 _25402_ (.A(_02182_),
    .B1(_01955_),
    .B2(_21665_),
    .ZN(_02183_));
 AOI21_X1 _25403_ (.A(_02176_),
    .B1(_02181_),
    .B2(_02183_),
    .ZN(_02184_));
 AOI21_X1 _25404_ (.A(_02179_),
    .B1(_02183_),
    .B2(_02174_),
    .ZN(_02185_));
 OAI21_X4 _25405_ (.A(_02179_),
    .B1(_02133_),
    .B2(_02139_),
    .ZN(_02186_));
 NOR2_X4 _25406_ (.A1(_02159_),
    .A2(_02186_),
    .ZN(_02187_));
 CLKBUF_X3 _25407_ (.A(_02161_),
    .Z(_02188_));
 NAND4_X2 _25408_ (.A1(_02188_),
    .A2(_02165_),
    .A3(_02089_),
    .A4(_02179_),
    .ZN(_02189_));
 OR4_X2 _25409_ (.A1(_01881_),
    .A2(_01846_),
    .A3(_01981_),
    .A4(_02001_),
    .ZN(_02190_));
 OAI21_X4 _25410_ (.A(_02121_),
    .B1(_02190_),
    .B2(_02027_),
    .ZN(_02191_));
 AOI21_X1 _25411_ (.A(_02191_),
    .B1(_02183_),
    .B2(_02161_),
    .ZN(_02192_));
 OAI21_X1 _25412_ (.A(_02192_),
    .B1(_02119_),
    .B2(_02090_),
    .ZN(_02193_));
 NAND2_X1 _25413_ (.A1(_02189_),
    .A2(_02193_),
    .ZN(_02194_));
 AOI21_X2 _25414_ (.A(_02185_),
    .B1(_02187_),
    .B2(_02194_),
    .ZN(_02195_));
 NAND2_X1 _25415_ (.A1(_02172_),
    .A2(_02145_),
    .ZN(_02196_));
 NOR2_X2 _25416_ (.A1(_02078_),
    .A2(_02196_),
    .ZN(_02197_));
 OR2_X1 _25417_ (.A1(_02195_),
    .A2(_02197_),
    .ZN(_02198_));
 INV_X1 _25418_ (.A(_02198_),
    .ZN(_02199_));
 AND2_X1 _25419_ (.A1(_02184_),
    .A2(_02199_),
    .ZN(_21674_));
 BUF_X4 _25420_ (.A(_01764_),
    .Z(_02200_));
 OR4_X1 _25421_ (.A1(\g_reduce0[4].adder.b[11] ),
    .A2(_01765_),
    .A3(_01766_),
    .A4(_01767_),
    .ZN(_02201_));
 CLKBUF_X3 _25422_ (.A(_02201_),
    .Z(_02202_));
 NAND2_X1 _25423_ (.A1(_01764_),
    .A2(_02202_),
    .ZN(_02203_));
 BUF_X4 _25424_ (.A(_02203_),
    .Z(_02204_));
 BUF_X1 _25425_ (.A(_21670_),
    .Z(_02205_));
 INV_X4 _25426_ (.A(_02159_),
    .ZN(_21696_));
 AND3_X1 _25427_ (.A1(_02205_),
    .A2(_21692_),
    .A3(_21696_),
    .ZN(_02206_));
 CLKBUF_X3 _25428_ (.A(_02145_),
    .Z(_02207_));
 OAI21_X1 _25429_ (.A(_02198_),
    .B1(_02206_),
    .B2(_02207_),
    .ZN(_02208_));
 MUX2_X1 _25430_ (.A(_02198_),
    .B(_02208_),
    .S(_02184_),
    .Z(_02209_));
 INV_X1 _25431_ (.A(_21677_),
    .ZN(_02210_));
 AOI21_X2 _25432_ (.A(_02030_),
    .B1(_02029_),
    .B2(_01905_),
    .ZN(_02211_));
 NOR3_X2 _25433_ (.A1(_02027_),
    .A2(_02026_),
    .A3(_02025_),
    .ZN(_02212_));
 NOR2_X2 _25434_ (.A1(_02211_),
    .A2(_02212_),
    .ZN(_02213_));
 NAND4_X2 _25435_ (.A1(_02188_),
    .A2(_02213_),
    .A3(_02099_),
    .A4(_02086_),
    .ZN(_02214_));
 OAI21_X1 _25436_ (.A(_02163_),
    .B1(_02165_),
    .B2(_02169_),
    .ZN(_02215_));
 NAND2_X1 _25437_ (.A1(_02214_),
    .A2(_02215_),
    .ZN(_02216_));
 AOI221_X2 _25438_ (.A(_02078_),
    .B1(_02187_),
    .B2(_02216_),
    .C1(_02085_),
    .C2(_02172_),
    .ZN(_02217_));
 OAI21_X1 _25439_ (.A(_02075_),
    .B1(_02125_),
    .B2(_02174_),
    .ZN(_02218_));
 NAND2_X1 _25440_ (.A1(_02207_),
    .A2(_02218_),
    .ZN(_02219_));
 NAND2_X1 _25441_ (.A1(_02188_),
    .A2(_02078_),
    .ZN(_02220_));
 NOR2_X2 _25442_ (.A1(_02090_),
    .A2(_02119_),
    .ZN(_02221_));
 CLKBUF_X3 _25443_ (.A(_02188_),
    .Z(_02222_));
 OAI221_X2 _25444_ (.A(_02214_),
    .B1(_02220_),
    .B2(_02221_),
    .C1(_02170_),
    .C2(_02222_),
    .ZN(_02223_));
 NAND2_X2 _25445_ (.A1(_02187_),
    .A2(_02223_),
    .ZN(_02224_));
 CLKBUF_X3 _25446_ (.A(_02140_),
    .Z(_02225_));
 AND2_X1 _25447_ (.A1(_02205_),
    .A2(_02225_),
    .ZN(_02226_));
 NAND2_X1 _25448_ (.A1(_02030_),
    .A2(_02099_),
    .ZN(_02227_));
 AOI21_X2 _25449_ (.A(_02227_),
    .B1(_02029_),
    .B2(_01904_),
    .ZN(_02228_));
 NOR4_X4 _25450_ (.A1(_02027_),
    .A2(_02026_),
    .A3(_02030_),
    .A4(_02083_),
    .ZN(_02229_));
 NOR3_X4 _25451_ (.A1(_02191_),
    .A2(_02228_),
    .A3(_02229_),
    .ZN(_02230_));
 AOI211_X2 _25452_ (.A(_02162_),
    .B(_02078_),
    .C1(_02230_),
    .C2(_02085_),
    .ZN(_02231_));
 NOR2_X1 _25453_ (.A1(_02162_),
    .A2(_02085_),
    .ZN(_02232_));
 NOR3_X1 _25454_ (.A1(_02183_),
    .A2(_02228_),
    .A3(_02229_),
    .ZN(_02233_));
 AND3_X1 _25455_ (.A1(_02028_),
    .A2(_02031_),
    .A3(_02089_),
    .ZN(_02234_));
 AOI21_X1 _25456_ (.A(_02233_),
    .B1(_02234_),
    .B2(_02165_),
    .ZN(_02235_));
 AOI221_X2 _25457_ (.A(_02231_),
    .B1(_02232_),
    .B2(_21669_),
    .C1(_02162_),
    .C2(_02235_),
    .ZN(_02236_));
 NOR2_X1 _25458_ (.A1(_02191_),
    .A2(_02140_),
    .ZN(_02237_));
 AOI21_X2 _25459_ (.A(_02226_),
    .B1(_02236_),
    .B2(_02237_),
    .ZN(_02238_));
 OAI22_X4 _25460_ (.A1(_02217_),
    .A2(_02219_),
    .B1(_02224_),
    .B2(_02238_),
    .ZN(_02239_));
 NOR3_X1 _25461_ (.A1(_02125_),
    .A2(_02075_),
    .A3(_02183_),
    .ZN(_02240_));
 NOR2_X1 _25462_ (.A1(_02196_),
    .A2(_02240_),
    .ZN(_02241_));
 NOR4_X4 _25463_ (.A1(_02176_),
    .A2(_02195_),
    .A3(_02197_),
    .A4(_02241_),
    .ZN(_02242_));
 NAND2_X1 _25464_ (.A1(_02239_),
    .A2(_02242_),
    .ZN(_02243_));
 MUX2_X1 _25465_ (.A(_02052_),
    .B(_02060_),
    .S(_02173_),
    .Z(_02244_));
 NAND2_X1 _25466_ (.A1(_02145_),
    .A2(_02244_),
    .ZN(_02245_));
 OAI21_X1 _25467_ (.A(_02245_),
    .B1(_02159_),
    .B2(_02145_),
    .ZN(_02246_));
 NAND2_X1 _25468_ (.A1(_21692_),
    .A2(_02245_),
    .ZN(_02247_));
 NOR2_X1 _25469_ (.A1(_02188_),
    .A2(_02125_),
    .ZN(_02248_));
 OAI21_X1 _25470_ (.A(_02248_),
    .B1(_02119_),
    .B2(_02090_),
    .ZN(_02249_));
 NAND2_X1 _25471_ (.A1(_02163_),
    .A2(_02085_),
    .ZN(_02250_));
 OAI21_X1 _25472_ (.A(_02083_),
    .B1(_02154_),
    .B2(_02156_),
    .ZN(_02251_));
 NAND2_X2 _25473_ (.A1(_02234_),
    .A2(_02251_),
    .ZN(_02252_));
 NOR2_X1 _25474_ (.A1(_02094_),
    .A2(_02099_),
    .ZN(_02253_));
 AOI21_X1 _25475_ (.A(_02065_),
    .B1(_02167_),
    .B2(_02168_),
    .ZN(_02254_));
 AOI21_X1 _25476_ (.A(_02094_),
    .B1(_02031_),
    .B2(_02028_),
    .ZN(_02255_));
 NOR3_X2 _25477_ (.A1(_02253_),
    .A2(_02254_),
    .A3(_02255_),
    .ZN(_02256_));
 OAI221_X2 _25478_ (.A(_02249_),
    .B1(_02250_),
    .B2(_02252_),
    .C1(_02256_),
    .C2(_02163_),
    .ZN(_02257_));
 OAI21_X1 _25479_ (.A(_02214_),
    .B1(_02220_),
    .B2(_02221_),
    .ZN(_02258_));
 NAND3_X1 _25480_ (.A1(_02225_),
    .A2(_02245_),
    .A3(_02215_),
    .ZN(_02259_));
 OAI221_X2 _25481_ (.A(_02246_),
    .B1(_02247_),
    .B2(_02257_),
    .C1(_02258_),
    .C2(_02259_),
    .ZN(_02260_));
 MUX2_X2 _25482_ (.A(_14111_),
    .B(_14107_),
    .S(_01984_),
    .Z(_02261_));
 NAND3_X2 _25483_ (.A1(_21672_),
    .A2(_02137_),
    .A3(_02138_),
    .ZN(_02262_));
 OAI21_X2 _25484_ (.A(_02120_),
    .B1(_02129_),
    .B2(_02132_),
    .ZN(_02263_));
 AOI21_X1 _25485_ (.A(_02261_),
    .B1(_02262_),
    .B2(_02263_),
    .ZN(_02264_));
 AOI21_X1 _25486_ (.A(_02183_),
    .B1(_02262_),
    .B2(_02263_),
    .ZN(_02265_));
 MUX2_X1 _25487_ (.A(_02264_),
    .B(_02265_),
    .S(_02221_),
    .Z(_02266_));
 NOR4_X2 _25488_ (.A1(_02222_),
    .A2(_02191_),
    .A3(_02144_),
    .A4(_02159_),
    .ZN(_02267_));
 NAND2_X1 _25489_ (.A1(_02188_),
    .A2(_02003_),
    .ZN(_02268_));
 NOR4_X2 _25490_ (.A1(_02165_),
    .A2(_02169_),
    .A3(_02133_),
    .A4(_02139_),
    .ZN(_02269_));
 NOR4_X1 _25491_ (.A1(_02145_),
    .A2(_02159_),
    .A3(_02268_),
    .A4(_02269_),
    .ZN(_02270_));
 NAND2_X2 _25492_ (.A1(_02068_),
    .A2(_02069_),
    .ZN(_02271_));
 OAI21_X2 _25493_ (.A(_02271_),
    .B1(_02090_),
    .B2(_02119_),
    .ZN(_02272_));
 OAI211_X2 _25494_ (.A(_02141_),
    .B(_02272_),
    .C1(_02075_),
    .C2(_02252_),
    .ZN(_02273_));
 MUX2_X1 _25495_ (.A(_02095_),
    .B(_02271_),
    .S(_02173_),
    .Z(_02274_));
 AOI222_X2 _25496_ (.A1(_02266_),
    .A2(_02267_),
    .B1(_02270_),
    .B2(_02273_),
    .C1(_02145_),
    .C2(_02274_),
    .ZN(_02275_));
 MUX2_X1 _25497_ (.A(_02094_),
    .B(_02065_),
    .S(_02173_),
    .Z(_02276_));
 NOR2_X1 _25498_ (.A1(_02179_),
    .A2(_02276_),
    .ZN(_02277_));
 NOR2_X1 _25499_ (.A1(_02162_),
    .A2(_02065_),
    .ZN(_02278_));
 OAI21_X1 _25500_ (.A(_02278_),
    .B1(_02230_),
    .B2(_02271_),
    .ZN(_02279_));
 OAI21_X2 _25501_ (.A(_02085_),
    .B1(_02078_),
    .B2(_02230_),
    .ZN(_02280_));
 MUX2_X1 _25502_ (.A(_02125_),
    .B(_02261_),
    .S(_02162_),
    .Z(_02281_));
 OAI221_X2 _25503_ (.A(_02279_),
    .B1(_02280_),
    .B2(_02188_),
    .C1(_21669_),
    .C2(_02281_),
    .ZN(_02282_));
 AOI211_X2 _25504_ (.A(_02144_),
    .B(_02159_),
    .C1(_02189_),
    .C2(_02193_),
    .ZN(_02283_));
 AOI221_X2 _25505_ (.A(_02277_),
    .B1(_02282_),
    .B2(_02187_),
    .C1(_02283_),
    .C2(_02225_),
    .ZN(_02284_));
 NOR3_X2 _25506_ (.A1(_02260_),
    .A2(_02275_),
    .A3(_02284_),
    .ZN(_02285_));
 MUX2_X1 _25507_ (.A(_02092_),
    .B(_02093_),
    .S(_02173_),
    .Z(_02286_));
 AOI22_X2 _25508_ (.A1(_02159_),
    .A2(_02171_),
    .B1(_02286_),
    .B2(_02145_),
    .ZN(_02287_));
 OAI211_X2 _25509_ (.A(_02222_),
    .B(_02272_),
    .C1(_02252_),
    .C2(_02075_),
    .ZN(_02288_));
 MUX2_X1 _25510_ (.A(_02078_),
    .B(_02086_),
    .S(_02221_),
    .Z(_02289_));
 OAI21_X1 _25511_ (.A(_02288_),
    .B1(_02289_),
    .B2(_02222_),
    .ZN(_02290_));
 NAND2_X1 _25512_ (.A1(_02225_),
    .A2(_02160_),
    .ZN(_02291_));
 OAI21_X1 _25513_ (.A(_02163_),
    .B1(_02191_),
    .B2(_02256_),
    .ZN(_02292_));
 NAND2_X1 _25514_ (.A1(_02028_),
    .A2(_02031_),
    .ZN(_02293_));
 AOI21_X1 _25515_ (.A(_02293_),
    .B1(_02091_),
    .B2(_02092_),
    .ZN(_02294_));
 OAI33_X1 _25516_ (.A1(_02084_),
    .A2(_02083_),
    .A3(_02145_),
    .B1(_02294_),
    .B2(_02191_),
    .B3(_02048_),
    .ZN(_02295_));
 OAI21_X1 _25517_ (.A(_02292_),
    .B1(_02295_),
    .B2(_02163_),
    .ZN(_02296_));
 NAND2_X1 _25518_ (.A1(_21692_),
    .A2(_02160_),
    .ZN(_02297_));
 OAI221_X2 _25519_ (.A(_02287_),
    .B1(_02290_),
    .B2(_02291_),
    .C1(_02296_),
    .C2(_02297_),
    .ZN(_02298_));
 MUX2_X1 _25520_ (.A(_02093_),
    .B(_02052_),
    .S(_02173_),
    .Z(_02299_));
 NOR2_X1 _25521_ (.A1(_02180_),
    .A2(_02299_),
    .ZN(_02300_));
 NAND2_X1 _25522_ (.A1(_02179_),
    .A2(_21696_),
    .ZN(_02301_));
 NOR2_X1 _25523_ (.A1(_02191_),
    .A2(_02234_),
    .ZN(_02302_));
 NAND2_X1 _25524_ (.A1(_02163_),
    .A2(_02165_),
    .ZN(_02303_));
 OAI22_X1 _25525_ (.A1(_02188_),
    .A2(_02140_),
    .B1(_02302_),
    .B2(_02303_),
    .ZN(_02304_));
 NOR3_X1 _25526_ (.A1(_02188_),
    .A2(_02183_),
    .A3(_21666_),
    .ZN(_02305_));
 OAI21_X1 _25527_ (.A(_02095_),
    .B1(_02271_),
    .B2(_02230_),
    .ZN(_02306_));
 OAI21_X1 _25528_ (.A(_02306_),
    .B1(_21669_),
    .B2(_02125_),
    .ZN(_02307_));
 OAI33_X1 _25529_ (.A1(_02301_),
    .A2(_02304_),
    .A3(_02305_),
    .B1(_02307_),
    .B2(_02186_),
    .B3(_02159_),
    .ZN(_02308_));
 OAI211_X2 _25530_ (.A(_02140_),
    .B(_02280_),
    .C1(_02261_),
    .C2(_21669_),
    .ZN(_02309_));
 NAND3_X1 _25531_ (.A1(_02094_),
    .A2(_21666_),
    .A3(_21692_),
    .ZN(_02310_));
 NAND3_X1 _25532_ (.A1(_02084_),
    .A2(_21669_),
    .A3(_21692_),
    .ZN(_02311_));
 NAND4_X1 _25533_ (.A1(_02222_),
    .A2(_02309_),
    .A3(_02310_),
    .A4(_02311_),
    .ZN(_02312_));
 AOI21_X1 _25534_ (.A(_21696_),
    .B1(_21692_),
    .B2(_02205_),
    .ZN(_02313_));
 AOI221_X2 _25535_ (.A(_02300_),
    .B1(_02308_),
    .B2(_02312_),
    .C1(_02313_),
    .C2(_02180_),
    .ZN(_02314_));
 NOR3_X1 _25536_ (.A1(_02211_),
    .A2(_02212_),
    .A3(_02048_),
    .ZN(_02315_));
 NAND3_X1 _25537_ (.A1(_02028_),
    .A2(_02031_),
    .A3(_02039_),
    .ZN(_02316_));
 AOI21_X1 _25538_ (.A(_02315_),
    .B1(_02316_),
    .B2(_02092_),
    .ZN(_02317_));
 NOR2_X1 _25539_ (.A1(_02163_),
    .A2(_02317_),
    .ZN(_02318_));
 MUX2_X1 _25540_ (.A(_02039_),
    .B(_02092_),
    .S(_02174_),
    .Z(_02319_));
 AOI22_X2 _25541_ (.A1(_02187_),
    .A2(_02318_),
    .B1(_02319_),
    .B2(_02207_),
    .ZN(_02320_));
 NOR2_X1 _25542_ (.A1(_02222_),
    .A2(_02225_),
    .ZN(_02321_));
 MUX2_X1 _25543_ (.A(_02052_),
    .B(_02060_),
    .S(_02221_),
    .Z(_02322_));
 AOI22_X2 _25544_ (.A1(_02225_),
    .A2(_02282_),
    .B1(_02321_),
    .B2(_02322_),
    .ZN(_02323_));
 NAND2_X1 _25545_ (.A1(_21669_),
    .A2(_02126_),
    .ZN(_02324_));
 MUX2_X1 _25546_ (.A(_02126_),
    .B(_02324_),
    .S(_21672_),
    .Z(_02325_));
 AOI21_X1 _25547_ (.A(_02135_),
    .B1(_02177_),
    .B2(_02178_),
    .ZN(_02326_));
 NAND4_X1 _25548_ (.A1(_02094_),
    .A2(_02065_),
    .A3(_02326_),
    .A4(_02194_),
    .ZN(_02327_));
 OAI221_X2 _25549_ (.A(_02320_),
    .B1(_02323_),
    .B2(_02301_),
    .C1(_02325_),
    .C2(_02327_),
    .ZN(_02328_));
 NAND4_X2 _25550_ (.A1(_02285_),
    .A2(_02298_),
    .A3(_02314_),
    .A4(_02328_),
    .ZN(_02329_));
 MUX2_X1 _25551_ (.A(_02293_),
    .B(_02039_),
    .S(_02174_),
    .Z(_02330_));
 NAND2_X1 _25552_ (.A1(_02207_),
    .A2(_02330_),
    .ZN(_02331_));
 NAND2_X1 _25553_ (.A1(_02003_),
    .A2(_02039_),
    .ZN(_02332_));
 AOI21_X1 _25554_ (.A(_02332_),
    .B1(_02041_),
    .B2(_02213_),
    .ZN(_02333_));
 AND2_X1 _25555_ (.A1(_02222_),
    .A2(_02333_),
    .ZN(_02334_));
 AOI21_X1 _25556_ (.A(_02334_),
    .B1(_02295_),
    .B2(_02163_),
    .ZN(_02335_));
 NOR2_X1 _25557_ (.A1(_21692_),
    .A2(_02159_),
    .ZN(_02336_));
 NOR2_X1 _25558_ (.A1(_02225_),
    .A2(_21696_),
    .ZN(_02337_));
 AOI22_X2 _25559_ (.A1(_02257_),
    .A2(_02336_),
    .B1(_02337_),
    .B2(_02223_),
    .ZN(_02338_));
 OAI221_X2 _25560_ (.A(_02331_),
    .B1(_02335_),
    .B2(_02186_),
    .C1(_02207_),
    .C2(_02338_),
    .ZN(_02339_));
 INV_X1 _25561_ (.A(_02339_),
    .ZN(_02340_));
 AOI221_X2 _25562_ (.A(_21696_),
    .B1(_02237_),
    .B2(_02236_),
    .C1(_02225_),
    .C2(_02205_),
    .ZN(_02341_));
 NAND2_X1 _25563_ (.A1(_02162_),
    .A2(_02048_),
    .ZN(_02342_));
 MUX2_X1 _25564_ (.A(_02162_),
    .B(_02342_),
    .S(_02039_),
    .Z(_02343_));
 OAI33_X1 _25565_ (.A1(_02188_),
    .A2(_02092_),
    .A3(_02315_),
    .B1(_02343_),
    .B2(_02212_),
    .B3(_02211_),
    .ZN(_02344_));
 NAND2_X1 _25566_ (.A1(_02095_),
    .A2(_02230_),
    .ZN(_02345_));
 NAND3_X2 _25567_ (.A1(_02162_),
    .A2(_02262_),
    .A3(_02263_),
    .ZN(_02346_));
 OAI221_X2 _25568_ (.A(_21696_),
    .B1(_02164_),
    .B2(_02344_),
    .C1(_02345_),
    .C2(_02346_),
    .ZN(_02347_));
 AOI221_X2 _25569_ (.A(_02346_),
    .B1(_02069_),
    .B2(_02068_),
    .C1(_02065_),
    .C2(_21669_),
    .ZN(_02348_));
 NOR2_X1 _25570_ (.A1(_02163_),
    .A2(_02141_),
    .ZN(_02349_));
 MUX2_X1 _25571_ (.A(_02052_),
    .B(_02060_),
    .S(_21666_),
    .Z(_02350_));
 AOI211_X2 _25572_ (.A(_02347_),
    .B(_02348_),
    .C1(_02349_),
    .C2(_02350_),
    .ZN(_02351_));
 NOR3_X2 _25573_ (.A1(_02191_),
    .A2(_02341_),
    .A3(_02351_),
    .ZN(_02352_));
 NAND2_X1 _25574_ (.A1(_02174_),
    .A2(_02213_),
    .ZN(_02353_));
 NOR3_X2 _25575_ (.A1(_02293_),
    .A2(_02341_),
    .A3(_02351_),
    .ZN(_02354_));
 NAND2_X1 _25576_ (.A1(_02172_),
    .A2(_02003_),
    .ZN(_02355_));
 OAI22_X1 _25577_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02354_),
    .B2(_02355_),
    .ZN(_02356_));
 NOR4_X2 _25578_ (.A1(_02243_),
    .A2(_02329_),
    .A3(_02340_),
    .A4(_02356_),
    .ZN(_02357_));
 NAND3_X1 _25579_ (.A1(_02222_),
    .A2(_02225_),
    .A3(_02295_),
    .ZN(_02358_));
 NOR2_X1 _25580_ (.A1(_02268_),
    .A2(_02269_),
    .ZN(_02359_));
 NOR2_X1 _25581_ (.A1(_02222_),
    .A2(_02164_),
    .ZN(_02360_));
 AOI22_X2 _25582_ (.A1(_02273_),
    .A2(_02359_),
    .B1(_02360_),
    .B2(_02289_),
    .ZN(_02361_));
 NOR3_X1 _25583_ (.A1(_02191_),
    .A2(_21692_),
    .A3(_02256_),
    .ZN(_02362_));
 AOI21_X1 _25584_ (.A(_02362_),
    .B1(_02333_),
    .B2(_21692_),
    .ZN(_02363_));
 OAI221_X2 _25585_ (.A(_02358_),
    .B1(_02361_),
    .B2(_21696_),
    .C1(_02222_),
    .C2(_02363_),
    .ZN(_02364_));
 AOI22_X4 _25586_ (.A1(_02174_),
    .A2(_02191_),
    .B1(_02180_),
    .B2(_02364_),
    .ZN(_02365_));
 XNOR2_X1 _25587_ (.A(_02357_),
    .B(_02365_),
    .ZN(_02366_));
 MUX2_X1 _25588_ (.A(_02209_),
    .B(_02210_),
    .S(_02366_),
    .Z(_02367_));
 NAND2_X4 _25589_ (.A1(_01764_),
    .A2(_01768_),
    .ZN(_02368_));
 OAI222_X1 _25590_ (.A1(_01812_),
    .A2(_02200_),
    .B1(_02204_),
    .B2(_02367_),
    .C1(_02368_),
    .C2(_01784_),
    .ZN(_00080_));
 OAI22_X4 _25591_ (.A1(\g_reduce0[4].adder.b[1] ),
    .A2(_02200_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[1] ),
    .ZN(_02369_));
 BUF_X4 _25592_ (.A(_02366_),
    .Z(_21680_));
 AND2_X1 _25593_ (.A1(_02187_),
    .A2(_02236_),
    .ZN(_02370_));
 MUX2_X1 _25594_ (.A(_02271_),
    .B(_02085_),
    .S(_02174_),
    .Z(_02371_));
 NAND2_X1 _25595_ (.A1(_02207_),
    .A2(_02371_),
    .ZN(_02372_));
 NAND2_X1 _25596_ (.A1(_02205_),
    .A2(_02225_),
    .ZN(_02373_));
 OAI21_X1 _25597_ (.A(_02372_),
    .B1(_02373_),
    .B2(_02301_),
    .ZN(_02374_));
 OAI21_X1 _25598_ (.A(_21676_),
    .B1(_02370_),
    .B2(_02374_),
    .ZN(_02375_));
 INV_X1 _25599_ (.A(_21676_),
    .ZN(_02376_));
 NAND2_X1 _25600_ (.A1(_02187_),
    .A2(_02236_),
    .ZN(_02377_));
 AOI22_X2 _25601_ (.A1(_02160_),
    .A2(_02226_),
    .B1(_02371_),
    .B2(_02207_),
    .ZN(_02378_));
 NAND3_X1 _25602_ (.A1(_02376_),
    .A2(_02377_),
    .A3(_02378_),
    .ZN(_02379_));
 AOI21_X1 _25603_ (.A(_02203_),
    .B1(_02375_),
    .B2(_02379_),
    .ZN(_02380_));
 AND2_X1 _25604_ (.A1(_21680_),
    .A2(_02380_),
    .ZN(_02381_));
 NOR3_X1 _25605_ (.A1(_21677_),
    .A2(_02204_),
    .A3(_21680_),
    .ZN(_02382_));
 NOR3_X1 _25606_ (.A1(_02369_),
    .A2(_02381_),
    .A3(_02382_),
    .ZN(_00087_));
 OAI22_X4 _25607_ (.A1(\g_reduce0[4].adder.b[2] ),
    .A2(_02200_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[2] ),
    .ZN(_02383_));
 AND2_X1 _25608_ (.A1(_02239_),
    .A2(_02242_),
    .ZN(_02384_));
 XNOR2_X1 _25609_ (.A(_02275_),
    .B(_02384_),
    .ZN(_02385_));
 NOR2_X1 _25610_ (.A1(_02204_),
    .A2(_02385_),
    .ZN(_02386_));
 MUX2_X1 _25611_ (.A(_02380_),
    .B(_02386_),
    .S(_21680_),
    .Z(_02387_));
 NOR2_X1 _25612_ (.A1(_02383_),
    .A2(_02387_),
    .ZN(_00088_));
 OAI22_X4 _25613_ (.A1(\g_reduce0[4].adder.b[3] ),
    .A2(_02200_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[3] ),
    .ZN(_02388_));
 OR2_X1 _25614_ (.A1(_02275_),
    .A2(_02375_),
    .ZN(_02389_));
 XOR2_X1 _25615_ (.A(_02284_),
    .B(_02389_),
    .Z(_02390_));
 NOR2_X1 _25616_ (.A1(_02204_),
    .A2(_02390_),
    .ZN(_02391_));
 MUX2_X1 _25617_ (.A(_02386_),
    .B(_02391_),
    .S(_21680_),
    .Z(_02392_));
 NOR2_X2 _25618_ (.A1(_02388_),
    .A2(_02392_),
    .ZN(_00089_));
 OAI22_X4 _25619_ (.A1(\g_reduce0[4].adder.b[4] ),
    .A2(_02200_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[4] ),
    .ZN(_02393_));
 NOR2_X1 _25620_ (.A1(_02275_),
    .A2(_02284_),
    .ZN(_02394_));
 NAND3_X1 _25621_ (.A1(_02394_),
    .A2(_02239_),
    .A3(_02242_),
    .ZN(_02395_));
 XOR2_X1 _25622_ (.A(_02260_),
    .B(_02395_),
    .Z(_02396_));
 OR2_X1 _25623_ (.A1(_02203_),
    .A2(_02396_),
    .ZN(_02397_));
 NAND2_X1 _25624_ (.A1(_21680_),
    .A2(_02397_),
    .ZN(_02398_));
 OR2_X1 _25625_ (.A1(_21680_),
    .A2(_02391_),
    .ZN(_02399_));
 AOI21_X2 _25626_ (.A(_02393_),
    .B1(_02398_),
    .B2(_02399_),
    .ZN(_00090_));
 NOR2_X1 _25627_ (.A1(_21680_),
    .A2(_02397_),
    .ZN(_02400_));
 AOI21_X2 _25628_ (.A(_02376_),
    .B1(_02377_),
    .B2(_02378_),
    .ZN(_02401_));
 NAND2_X1 _25629_ (.A1(_02285_),
    .A2(_02401_),
    .ZN(_02402_));
 XNOR2_X1 _25630_ (.A(_02314_),
    .B(_02402_),
    .ZN(_02403_));
 NOR2_X1 _25631_ (.A1(_02204_),
    .A2(_02403_),
    .ZN(_02404_));
 NOR4_X4 _25632_ (.A1(\g_reduce0[4].adder.a[11] ),
    .A2(_01761_),
    .A3(\g_reduce0[4].adder.a[14] ),
    .A4(_01762_),
    .ZN(_02405_));
 NAND2_X1 _25633_ (.A1(\g_reduce0[4].adder.b[5] ),
    .A2(_02405_),
    .ZN(_02406_));
 OAI21_X1 _25634_ (.A(_01764_),
    .B1(_02202_),
    .B2(\g_reduce0[4].adder.a[5] ),
    .ZN(_02407_));
 AOI221_X1 _25635_ (.A(_02400_),
    .B1(_02404_),
    .B2(_21680_),
    .C1(_02406_),
    .C2(_02407_),
    .ZN(_00091_));
 OAI22_X2 _25636_ (.A1(\g_reduce0[4].adder.b[6] ),
    .A2(_01764_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[6] ),
    .ZN(_02408_));
 NOR2_X1 _25637_ (.A1(_02243_),
    .A2(_02329_),
    .ZN(_02409_));
 NOR2_X2 _25638_ (.A1(_02340_),
    .A2(_02356_),
    .ZN(_02410_));
 NAND2_X1 _25639_ (.A1(_02409_),
    .A2(_02410_),
    .ZN(_02411_));
 BUF_X2 _25640_ (.A(_02365_),
    .Z(_02412_));
 AND2_X1 _25641_ (.A1(_02412_),
    .A2(_02403_),
    .ZN(_02413_));
 AOI21_X1 _25642_ (.A(_02204_),
    .B1(_02411_),
    .B2(_02413_),
    .ZN(_02414_));
 NAND4_X2 _25643_ (.A1(_02285_),
    .A2(_02314_),
    .A3(_02239_),
    .A4(_02242_),
    .ZN(_02415_));
 XNOR2_X2 _25644_ (.A(_02298_),
    .B(_02415_),
    .ZN(_02416_));
 AOI21_X1 _25645_ (.A(_02416_),
    .B1(_02403_),
    .B2(_02357_),
    .ZN(_02417_));
 OR2_X1 _25646_ (.A1(_02412_),
    .A2(_02417_),
    .ZN(_02418_));
 AOI21_X2 _25647_ (.A(_02408_),
    .B1(_02414_),
    .B2(_02418_),
    .ZN(_00092_));
 OAI22_X2 _25648_ (.A1(\g_reduce0[4].adder.b[7] ),
    .A2(_02200_),
    .B1(_02368_),
    .B2(\g_reduce0[4].adder.a[7] ),
    .ZN(_02419_));
 AND4_X1 _25649_ (.A1(_02285_),
    .A2(_02298_),
    .A3(_02314_),
    .A4(_02401_),
    .ZN(_02420_));
 XOR2_X2 _25650_ (.A(_02328_),
    .B(_02420_),
    .Z(_02421_));
 AOI221_X2 _25651_ (.A(_02204_),
    .B1(_02412_),
    .B2(_02416_),
    .C1(_02421_),
    .C2(_21680_),
    .ZN(_02422_));
 NOR2_X2 _25652_ (.A1(_02419_),
    .A2(_02422_),
    .ZN(_00093_));
 NAND2_X2 _25653_ (.A1(\g_reduce0[4].adder.b[8] ),
    .A2(_02405_),
    .ZN(_02423_));
 NAND2_X1 _25654_ (.A1(_02202_),
    .A2(_02412_),
    .ZN(_02424_));
 OAI221_X2 _25655_ (.A(_01764_),
    .B1(_02411_),
    .B2(_02424_),
    .C1(_02202_),
    .C2(\g_reduce0[4].adder.a[8] ),
    .ZN(_02425_));
 XNOR2_X1 _25656_ (.A(_02409_),
    .B(_02339_),
    .ZN(_02426_));
 OR2_X1 _25657_ (.A1(_02412_),
    .A2(_02426_),
    .ZN(_02427_));
 OR2_X1 _25658_ (.A1(_02204_),
    .A2(_02412_),
    .ZN(_02428_));
 OAI22_X4 _25659_ (.A1(_02410_),
    .A2(_02428_),
    .B1(_02421_),
    .B2(_02204_),
    .ZN(_02429_));
 AOI22_X4 _25660_ (.A1(_02423_),
    .A2(_02425_),
    .B1(_02427_),
    .B2(_02429_),
    .ZN(_00094_));
 NOR4_X1 _25661_ (.A1(_02384_),
    .A2(_02356_),
    .A3(_02365_),
    .A4(_02401_),
    .ZN(_02430_));
 NOR3_X1 _25662_ (.A1(_02340_),
    .A2(_02412_),
    .A3(_02375_),
    .ZN(_02431_));
 AOI21_X1 _25663_ (.A(_02430_),
    .B1(_02431_),
    .B2(_02356_),
    .ZN(_02432_));
 MUX2_X1 _25664_ (.A(_02356_),
    .B(_02340_),
    .S(_02365_),
    .Z(_02433_));
 MUX2_X1 _25665_ (.A(_02432_),
    .B(_02433_),
    .S(_02329_),
    .Z(_02434_));
 OAI21_X1 _25666_ (.A(_02339_),
    .B1(_02356_),
    .B2(_02401_),
    .ZN(_02435_));
 AND3_X1 _25667_ (.A1(_02409_),
    .A2(_02412_),
    .A3(_02435_),
    .ZN(_02436_));
 NOR3_X2 _25668_ (.A1(_02339_),
    .A2(_02356_),
    .A3(_02412_),
    .ZN(_02437_));
 AND3_X1 _25669_ (.A1(_02243_),
    .A2(_02339_),
    .A3(_02412_),
    .ZN(_02438_));
 NOR4_X4 _25670_ (.A1(_02204_),
    .A2(_02436_),
    .A3(_02437_),
    .A4(_02438_),
    .ZN(_02439_));
 NAND2_X1 _25671_ (.A1(\g_reduce0[4].adder.b[9] ),
    .A2(_02405_),
    .ZN(_02440_));
 OAI21_X2 _25672_ (.A(_01764_),
    .B1(_02202_),
    .B2(\g_reduce0[4].adder.a[9] ),
    .ZN(_02441_));
 AOI22_X4 _25673_ (.A1(_02434_),
    .A2(_02439_),
    .B1(_02440_),
    .B2(_02441_),
    .ZN(_00095_));
 INV_X1 _25674_ (.A(_21684_),
    .ZN(_21678_));
 MUX2_X1 _25675_ (.A(\g_reduce0[4].adder.a[10] ),
    .B(_21683_),
    .S(_02202_),
    .Z(_02442_));
 MUX2_X2 _25676_ (.A(\g_reduce0[4].adder.b[10] ),
    .B(_02442_),
    .S(_02200_),
    .Z(_00081_));
 MUX2_X1 _25677_ (.A(\g_reduce0[4].adder.a[11] ),
    .B(_21691_),
    .S(_02202_),
    .Z(_02443_));
 MUX2_X2 _25678_ (.A(\g_reduce0[4].adder.b[11] ),
    .B(_02443_),
    .S(_02200_),
    .Z(_00082_));
 MUX2_X2 _25679_ (.A(_21559_),
    .B(_00528_),
    .S(_01821_),
    .Z(_02444_));
 NAND2_X1 _25680_ (.A1(_02172_),
    .A2(_21685_),
    .ZN(_02445_));
 XOR2_X1 _25681_ (.A(_02444_),
    .B(_02445_),
    .Z(_02446_));
 XOR2_X1 _25682_ (.A(_14115_),
    .B(_21695_),
    .Z(_02447_));
 MUX2_X1 _25683_ (.A(_02446_),
    .B(_02447_),
    .S(_02180_),
    .Z(_02448_));
 XOR2_X1 _25684_ (.A(_21690_),
    .B(_02448_),
    .Z(_02449_));
 MUX2_X1 _25685_ (.A(_01761_),
    .B(_02449_),
    .S(_02202_),
    .Z(_02450_));
 MUX2_X2 _25686_ (.A(_01765_),
    .B(_02450_),
    .S(_02200_),
    .Z(_00083_));
 INV_X1 _25687_ (.A(_14117_),
    .ZN(_14114_));
 MUX2_X1 _25688_ (.A(_21556_),
    .B(_00531_),
    .S(_01821_),
    .Z(_02451_));
 MUX2_X1 _25689_ (.A(_21562_),
    .B(_00523_),
    .S(_01821_),
    .Z(_02452_));
 NAND2_X1 _25690_ (.A1(_02172_),
    .A2(_21684_),
    .ZN(_02453_));
 NOR3_X1 _25691_ (.A1(_02444_),
    .A2(_02452_),
    .A3(_02453_),
    .ZN(_02454_));
 XNOR2_X1 _25692_ (.A(_02451_),
    .B(_02454_),
    .ZN(_02455_));
 INV_X1 _25693_ (.A(_21687_),
    .ZN(_02456_));
 INV_X1 _25694_ (.A(_21688_),
    .ZN(_02457_));
 OAI21_X1 _25695_ (.A(_02456_),
    .B1(_02457_),
    .B2(_14117_),
    .ZN(_02458_));
 AOI21_X1 _25696_ (.A(_21694_),
    .B1(_02458_),
    .B2(_21695_),
    .ZN(_02459_));
 XNOR2_X1 _25697_ (.A(_21699_),
    .B(_02459_),
    .ZN(_02460_));
 MUX2_X1 _25698_ (.A(_02455_),
    .B(_02460_),
    .S(_02180_),
    .Z(_02461_));
 NAND2_X1 _25699_ (.A1(_02172_),
    .A2(_21686_),
    .ZN(_02462_));
 OAI21_X1 _25700_ (.A(_02462_),
    .B1(_02452_),
    .B2(_02172_),
    .ZN(_02463_));
 MUX2_X1 _25701_ (.A(_14116_),
    .B(_02463_),
    .S(_02207_),
    .Z(_21689_));
 NAND3_X1 _25702_ (.A1(_21682_),
    .A2(_02448_),
    .A3(_21689_),
    .ZN(_02464_));
 XNOR2_X1 _25703_ (.A(_02461_),
    .B(_02464_),
    .ZN(_02465_));
 MUX2_X1 _25704_ (.A(\g_reduce0[4].adder.a[13] ),
    .B(_02465_),
    .S(_02202_),
    .Z(_02466_));
 MUX2_X2 _25705_ (.A(\g_reduce0[4].adder.b[13] ),
    .B(_02466_),
    .S(_02200_),
    .Z(_00084_));
 OR2_X1 _25706_ (.A1(_01766_),
    .A2(_01805_),
    .ZN(_02467_));
 NAND2_X1 _25707_ (.A1(\g_reduce0[4].adder.a[14] ),
    .A2(_02467_),
    .ZN(_02468_));
 NOR4_X1 _25708_ (.A1(_02180_),
    .A2(_02444_),
    .A3(_02445_),
    .A4(_02451_),
    .ZN(_02469_));
 AOI21_X1 _25709_ (.A(_21694_),
    .B1(_21695_),
    .B2(_14115_),
    .ZN(_02470_));
 INV_X1 _25710_ (.A(_02470_),
    .ZN(_02471_));
 AOI21_X1 _25711_ (.A(_21698_),
    .B1(_02471_),
    .B2(_21699_),
    .ZN(_02472_));
 AOI21_X1 _25712_ (.A(_02469_),
    .B1(_02472_),
    .B2(_02180_),
    .ZN(_02473_));
 NAND3_X1 _25713_ (.A1(_21690_),
    .A2(_02448_),
    .A3(_02461_),
    .ZN(_02474_));
 XOR2_X2 _25714_ (.A(_02473_),
    .B(_02474_),
    .Z(_02475_));
 MUX2_X1 _25715_ (.A(_02467_),
    .B(_02468_),
    .S(_02475_),
    .Z(_02476_));
 OAI22_X1 _25716_ (.A1(_01766_),
    .A2(_01764_),
    .B1(_01768_),
    .B2(_02476_),
    .ZN(_02477_));
 NOR2_X1 _25717_ (.A1(\g_reduce0[4].adder.a[14] ),
    .A2(_02405_),
    .ZN(_02478_));
 NAND3_X1 _25718_ (.A1(_01766_),
    .A2(_01849_),
    .A3(_02475_),
    .ZN(_02479_));
 OR2_X1 _25719_ (.A1(_01849_),
    .A2(_02475_),
    .ZN(_02480_));
 NAND3_X1 _25720_ (.A1(_02202_),
    .A2(_02479_),
    .A3(_02480_),
    .ZN(_02481_));
 AOI21_X1 _25721_ (.A(_02477_),
    .B1(_02478_),
    .B2(_02481_),
    .ZN(_00085_));
 BUF_X2 _25722_ (.A(\g_reduce0[6].adder.a[11] ),
    .Z(_02482_));
 BUF_X2 _25723_ (.A(\g_reduce0[6].adder.a[12] ),
    .Z(_02483_));
 BUF_X2 _25724_ (.A(\g_reduce0[6].adder.a[14] ),
    .Z(_02484_));
 OR2_X1 _25725_ (.A1(\g_reduce0[6].adder.a[10] ),
    .A2(\g_reduce0[6].adder.a[13] ),
    .ZN(_02485_));
 OR4_X2 _25726_ (.A1(_02482_),
    .A2(_02483_),
    .A3(_02484_),
    .A4(_02485_),
    .ZN(_02486_));
 CLKBUF_X2 _25727_ (.A(\g_reduce0[6].adder.b[11] ),
    .Z(_02487_));
 CLKBUF_X2 _25728_ (.A(\g_reduce0[6].adder.b[12] ),
    .Z(_02488_));
 BUF_X2 _25729_ (.A(\g_reduce0[6].adder.b[14] ),
    .Z(_02489_));
 OR2_X1 _25730_ (.A1(\g_reduce0[6].adder.b[10] ),
    .A2(\g_reduce0[6].adder.b[13] ),
    .ZN(_02490_));
 NOR4_X4 _25731_ (.A1(_02487_),
    .A2(_02488_),
    .A3(_02489_),
    .A4(_02490_),
    .ZN(_02491_));
 INV_X1 _25732_ (.A(_21746_),
    .ZN(_02492_));
 BUF_X4 _25733_ (.A(_21702_),
    .Z(_02493_));
 AOI21_X2 _25734_ (.A(_21701_),
    .B1(_21704_),
    .B2(_02493_),
    .ZN(_02494_));
 BUF_X2 _25735_ (.A(_21747_),
    .Z(_02495_));
 INV_X1 _25736_ (.A(_02495_),
    .ZN(_02496_));
 OAI21_X2 _25737_ (.A(_02492_),
    .B1(_02494_),
    .B2(_02496_),
    .ZN(_02497_));
 BUF_X4 _25738_ (.A(_21705_),
    .Z(_02498_));
 INV_X2 _25739_ (.A(_02498_),
    .ZN(_02499_));
 NAND2_X1 _25740_ (.A1(_02495_),
    .A2(_02493_),
    .ZN(_02500_));
 NOR2_X2 _25741_ (.A1(_02499_),
    .A2(_02500_),
    .ZN(_02501_));
 INV_X1 _25742_ (.A(_21707_),
    .ZN(_02502_));
 INV_X1 _25743_ (.A(_21708_),
    .ZN(_02503_));
 OAI21_X2 _25744_ (.A(_02502_),
    .B1(_21740_),
    .B2(_02503_),
    .ZN(_02504_));
 AOI21_X4 _25745_ (.A(_02497_),
    .B1(_02501_),
    .B2(_02504_),
    .ZN(_02505_));
 BUF_X2 _25746_ (.A(_21741_),
    .Z(_02506_));
 AND2_X1 _25747_ (.A1(_02495_),
    .A2(_02493_),
    .ZN(_02507_));
 AND2_X2 _25748_ (.A1(_02498_),
    .A2(_21708_),
    .ZN(_02508_));
 AND3_X1 _25749_ (.A1(_02506_),
    .A2(_02507_),
    .A3(_02508_),
    .ZN(_02509_));
 INV_X1 _25750_ (.A(_21710_),
    .ZN(_02510_));
 AOI211_X2 _25751_ (.A(_21713_),
    .B(_21716_),
    .C1(_21719_),
    .C2(_21717_),
    .ZN(_02511_));
 OAI21_X1 _25752_ (.A(_21711_),
    .B1(_21714_),
    .B2(_21713_),
    .ZN(_02512_));
 OAI21_X1 _25753_ (.A(_02510_),
    .B1(_02511_),
    .B2(_02512_),
    .ZN(_02513_));
 AOI21_X1 _25754_ (.A(_21722_),
    .B1(_21725_),
    .B2(_21723_),
    .ZN(_02514_));
 AOI21_X1 _25755_ (.A(_21728_),
    .B1(_21729_),
    .B2(_21731_),
    .ZN(_02515_));
 NAND2_X1 _25756_ (.A1(_21723_),
    .A2(_21726_),
    .ZN(_02516_));
 OAI21_X1 _25757_ (.A(_02514_),
    .B1(_02515_),
    .B2(_02516_),
    .ZN(_02517_));
 NAND4_X4 _25758_ (.A1(_21711_),
    .A2(_21714_),
    .A3(_21717_),
    .A4(_21720_),
    .ZN(_02518_));
 INV_X1 _25759_ (.A(_02518_),
    .ZN(_02519_));
 NAND4_X2 _25760_ (.A1(_21723_),
    .A2(_21726_),
    .A3(_21729_),
    .A4(_21732_),
    .ZN(_02520_));
 NOR2_X1 _25761_ (.A1(_02518_),
    .A2(_02520_),
    .ZN(_02521_));
 INV_X1 _25762_ (.A(_21734_),
    .ZN(_02522_));
 INV_X1 _25763_ (.A(_21735_),
    .ZN(_02523_));
 OAI21_X1 _25764_ (.A(_02522_),
    .B1(_21737_),
    .B2(_02523_),
    .ZN(_02524_));
 AOI221_X2 _25765_ (.A(_02513_),
    .B1(_02517_),
    .B2(_02519_),
    .C1(_02521_),
    .C2(_02524_),
    .ZN(_02525_));
 BUF_X4 _25766_ (.A(_02525_),
    .Z(_02526_));
 NAND3_X4 _25767_ (.A1(_02506_),
    .A2(_02507_),
    .A3(_02508_),
    .ZN(_02527_));
 NAND2_X1 _25768_ (.A1(_21735_),
    .A2(_21738_),
    .ZN(_02528_));
 NOR3_X4 _25769_ (.A1(_02518_),
    .A2(_02520_),
    .A3(_02528_),
    .ZN(_02529_));
 OR2_X2 _25770_ (.A1(_02527_),
    .A2(_02529_),
    .ZN(_02530_));
 OAI22_X4 _25771_ (.A1(_02505_),
    .A2(_02509_),
    .B1(_02526_),
    .B2(_02530_),
    .ZN(_02531_));
 BUF_X4 _25772_ (.A(_02531_),
    .Z(_02532_));
 CLKBUF_X3 _25773_ (.A(_02532_),
    .Z(_02533_));
 OAI21_X1 _25774_ (.A(_02486_),
    .B1(_02491_),
    .B2(_02533_),
    .ZN(_02534_));
 MUX2_X1 _25775_ (.A(\g_reduce0[6].adder.a[15] ),
    .B(\g_reduce0[6].adder.b[15] ),
    .S(_02534_),
    .Z(_00102_));
 MUX2_X2 _25776_ (.A(_00534_),
    .B(_21739_),
    .S(_02532_),
    .Z(_21825_));
 OR2_X1 _25777_ (.A1(_02488_),
    .A2(_00542_),
    .ZN(_02535_));
 NOR3_X1 _25778_ (.A1(_02526_),
    .A2(_02530_),
    .A3(_02535_),
    .ZN(_02536_));
 OR2_X1 _25779_ (.A1(_02483_),
    .A2(_21703_),
    .ZN(_02537_));
 NOR2_X1 _25780_ (.A1(_02527_),
    .A2(_02537_),
    .ZN(_02538_));
 OR2_X1 _25781_ (.A1(_02526_),
    .A2(_02529_),
    .ZN(_02539_));
 NOR2_X1 _25782_ (.A1(_02483_),
    .A2(_21703_),
    .ZN(_02540_));
 NOR2_X1 _25783_ (.A1(_02488_),
    .A2(_00542_),
    .ZN(_02541_));
 INV_X1 _25784_ (.A(_21740_),
    .ZN(_02542_));
 AOI21_X1 _25785_ (.A(_21707_),
    .B1(_02542_),
    .B2(_21708_),
    .ZN(_02543_));
 NAND2_X1 _25786_ (.A1(_02498_),
    .A2(_02507_),
    .ZN(_02544_));
 OAI221_X2 _25787_ (.A(_02492_),
    .B1(_02543_),
    .B2(_02544_),
    .C1(_02494_),
    .C2(_02496_),
    .ZN(_02545_));
 MUX2_X1 _25788_ (.A(_02540_),
    .B(_02541_),
    .S(_02545_),
    .Z(_02546_));
 AOI221_X2 _25789_ (.A(_02536_),
    .B1(_02538_),
    .B2(_02539_),
    .C1(_02527_),
    .C2(_02546_),
    .ZN(_02547_));
 OR2_X1 _25790_ (.A1(_02526_),
    .A2(_02530_),
    .ZN(_02548_));
 OR2_X1 _25791_ (.A1(\g_reduce0[6].adder.a[13] ),
    .A2(_21700_),
    .ZN(_02549_));
 AOI21_X1 _25792_ (.A(_02549_),
    .B1(_02527_),
    .B2(_02545_),
    .ZN(_02550_));
 NOR2_X1 _25793_ (.A1(\g_reduce0[6].adder.b[13] ),
    .A2(_00545_),
    .ZN(_02551_));
 AOI221_X2 _25794_ (.A(_02495_),
    .B1(_02548_),
    .B2(_02550_),
    .C1(_02551_),
    .C2(_02532_),
    .ZN(_02552_));
 INV_X1 _25795_ (.A(_21743_),
    .ZN(_02553_));
 NOR3_X1 _25796_ (.A1(_02482_),
    .A2(_21706_),
    .A3(_02527_),
    .ZN(_02554_));
 OAI21_X2 _25797_ (.A(_02554_),
    .B1(_02529_),
    .B2(_02526_),
    .ZN(_02555_));
 OR4_X2 _25798_ (.A1(_02487_),
    .A2(_00537_),
    .A3(_02526_),
    .A4(_02530_),
    .ZN(_02556_));
 OR3_X1 _25799_ (.A1(_02487_),
    .A2(_00537_),
    .A3(_02509_),
    .ZN(_02557_));
 OR3_X1 _25800_ (.A1(_02482_),
    .A2(_21706_),
    .A3(_02509_),
    .ZN(_02558_));
 MUX2_X2 _25801_ (.A(_02557_),
    .B(_02558_),
    .S(_02505_),
    .Z(_02559_));
 AND4_X2 _25802_ (.A1(_02553_),
    .A2(_02555_),
    .A3(_02556_),
    .A4(_02559_),
    .ZN(_02560_));
 OAI211_X4 _25803_ (.A(_02547_),
    .B(_02552_),
    .C1(_02499_),
    .C2(_02560_),
    .ZN(_02561_));
 NAND4_X4 _25804_ (.A1(_02553_),
    .A2(_02555_),
    .A3(_02556_),
    .A4(_02559_),
    .ZN(_02562_));
 OAI21_X1 _25805_ (.A(_02538_),
    .B1(_02529_),
    .B2(_02526_),
    .ZN(_02563_));
 MUX2_X1 _25806_ (.A(_02537_),
    .B(_02535_),
    .S(_02545_),
    .Z(_02564_));
 OAI221_X2 _25807_ (.A(_02563_),
    .B1(_02535_),
    .B2(_02548_),
    .C1(_02564_),
    .C2(_02509_),
    .ZN(_02565_));
 AOI22_X4 _25808_ (.A1(_02501_),
    .A2(_02562_),
    .B1(_02565_),
    .B2(_02507_),
    .ZN(_02566_));
 INV_X2 _25809_ (.A(_02493_),
    .ZN(_02567_));
 NAND2_X1 _25810_ (.A1(_02496_),
    .A2(_02567_),
    .ZN(_02568_));
 NOR2_X1 _25811_ (.A1(\g_reduce0[6].adder.a[13] ),
    .A2(_21700_),
    .ZN(_02569_));
 MUX2_X1 _25812_ (.A(_02569_),
    .B(_02551_),
    .S(_02532_),
    .Z(_02570_));
 MUX2_X2 _25813_ (.A(_02568_),
    .B(_02496_),
    .S(_02570_),
    .Z(_02571_));
 NAND3_X4 _25814_ (.A1(_02561_),
    .A2(_02566_),
    .A3(_02571_),
    .ZN(_02572_));
 INV_X1 _25815_ (.A(_21739_),
    .ZN(_02573_));
 NOR4_X1 _25816_ (.A1(_00534_),
    .A2(_02573_),
    .A3(_02527_),
    .A4(_02529_),
    .ZN(_02574_));
 AND2_X1 _25817_ (.A1(_00534_),
    .A2(_02573_),
    .ZN(_02575_));
 AND2_X1 _25818_ (.A1(_02509_),
    .A2(_02575_),
    .ZN(_02576_));
 MUX2_X1 _25819_ (.A(_02574_),
    .B(_02576_),
    .S(_02526_),
    .Z(_02577_));
 MUX2_X1 _25820_ (.A(_02505_),
    .B(_02529_),
    .S(_02509_),
    .Z(_02578_));
 NOR2_X1 _25821_ (.A1(_00534_),
    .A2(_02573_),
    .ZN(_02579_));
 NOR2_X1 _25822_ (.A1(_02505_),
    .A2(_02509_),
    .ZN(_02580_));
 AOI221_X1 _25823_ (.A(_02577_),
    .B1(_02578_),
    .B2(_02575_),
    .C1(_02579_),
    .C2(_02580_),
    .ZN(_21742_));
 NAND3_X1 _25824_ (.A1(_02555_),
    .A2(_02556_),
    .A3(_02559_),
    .ZN(_02581_));
 AOI221_X2 _25825_ (.A(_02565_),
    .B1(_21742_),
    .B2(_02508_),
    .C1(_02581_),
    .C2(_02498_),
    .ZN(_02582_));
 BUF_X4 _25826_ (.A(_02582_),
    .Z(_02583_));
 XNOR2_X2 _25827_ (.A(_02493_),
    .B(_02583_),
    .ZN(_02584_));
 MUX2_X1 _25828_ (.A(_00536_),
    .B(_21730_),
    .S(_02533_),
    .Z(_02585_));
 MUX2_X1 _25829_ (.A(_21736_),
    .B(_00533_),
    .S(_02533_),
    .Z(_02586_));
 BUF_X1 _25830_ (.A(_21744_),
    .Z(_02587_));
 BUF_X1 _25831_ (.A(_02587_),
    .Z(_02588_));
 INV_X1 _25832_ (.A(_02588_),
    .ZN(_02589_));
 MUX2_X1 _25833_ (.A(_02585_),
    .B(_02586_),
    .S(_02589_),
    .Z(_02590_));
 MUX2_X1 _25834_ (.A(_00535_),
    .B(_21727_),
    .S(_02533_),
    .Z(_02591_));
 NOR2_X1 _25835_ (.A1(_02589_),
    .A2(_02591_),
    .ZN(_02592_));
 INV_X1 _25836_ (.A(_00532_),
    .ZN(_02593_));
 INV_X1 _25837_ (.A(_21733_),
    .ZN(_02594_));
 MUX2_X1 _25838_ (.A(_02593_),
    .B(_02594_),
    .S(_02531_),
    .Z(_02595_));
 AOI21_X1 _25839_ (.A(_02592_),
    .B1(_02595_),
    .B2(_02589_),
    .ZN(_02596_));
 CLKBUF_X3 _25840_ (.A(_02506_),
    .Z(_02597_));
 INV_X2 _25841_ (.A(_02597_),
    .ZN(_02598_));
 MUX2_X1 _25842_ (.A(_02590_),
    .B(_02596_),
    .S(_02598_),
    .Z(_02599_));
 MUX2_X1 _25843_ (.A(_00538_),
    .B(_21721_),
    .S(_02533_),
    .Z(_02600_));
 MUX2_X1 _25844_ (.A(_00540_),
    .B(_21715_),
    .S(_02532_),
    .Z(_02601_));
 MUX2_X1 _25845_ (.A(_02600_),
    .B(_02601_),
    .S(_02588_),
    .Z(_02602_));
 MUX2_X1 _25846_ (.A(_00539_),
    .B(_21724_),
    .S(_02533_),
    .Z(_02603_));
 MUX2_X1 _25847_ (.A(_00541_),
    .B(_21718_),
    .S(_02533_),
    .Z(_02604_));
 MUX2_X1 _25848_ (.A(_02603_),
    .B(_02604_),
    .S(_02588_),
    .Z(_02605_));
 MUX2_X1 _25849_ (.A(_02602_),
    .B(_02605_),
    .S(_02597_),
    .Z(_02606_));
 XNOR2_X1 _25850_ (.A(_02498_),
    .B(_02560_),
    .ZN(_02607_));
 CLKBUF_X3 _25851_ (.A(_02607_),
    .Z(_02608_));
 MUX2_X1 _25852_ (.A(_02599_),
    .B(_02606_),
    .S(_02608_),
    .Z(_02609_));
 XNOR2_X2 _25853_ (.A(_02499_),
    .B(_02560_),
    .ZN(_02610_));
 CLKBUF_X3 _25854_ (.A(_02610_),
    .Z(_02611_));
 NAND2_X1 _25855_ (.A1(_02611_),
    .A2(_02584_),
    .ZN(_02612_));
 NAND2_X1 _25856_ (.A1(_02598_),
    .A2(_02587_),
    .ZN(_02613_));
 MUX2_X1 _25857_ (.A(_00543_),
    .B(_21709_),
    .S(_02532_),
    .Z(_02614_));
 OR2_X1 _25858_ (.A1(_02597_),
    .A2(_02614_),
    .ZN(_02615_));
 MUX2_X1 _25859_ (.A(_00544_),
    .B(_21712_),
    .S(_02532_),
    .Z(_02616_));
 OAI21_X1 _25860_ (.A(_02615_),
    .B1(_02616_),
    .B2(_02598_),
    .ZN(_02617_));
 OAI21_X1 _25861_ (.A(_02613_),
    .B1(_02617_),
    .B2(_02588_),
    .ZN(_02618_));
 OAI22_X1 _25862_ (.A1(_02584_),
    .A2(_02609_),
    .B1(_02612_),
    .B2(_02618_),
    .ZN(_02619_));
 NAND2_X1 _25863_ (.A1(_02572_),
    .A2(_02619_),
    .ZN(_21811_));
 INV_X1 _25864_ (.A(_21811_),
    .ZN(_21808_));
 XNOR2_X2 _25865_ (.A(_02567_),
    .B(_02583_),
    .ZN(_02620_));
 MUX2_X1 _25866_ (.A(_02585_),
    .B(_02603_),
    .S(_02588_),
    .Z(_02621_));
 MUX2_X1 _25867_ (.A(_02596_),
    .B(_02621_),
    .S(_02598_),
    .Z(_02622_));
 NAND2_X1 _25868_ (.A1(_02620_),
    .A2(_02622_),
    .ZN(_02623_));
 AOI21_X2 _25869_ (.A(_02588_),
    .B1(_02614_),
    .B2(_02597_),
    .ZN(_02624_));
 OAI21_X1 _25870_ (.A(_02623_),
    .B1(_02624_),
    .B2(_02620_),
    .ZN(_02625_));
 MUX2_X1 _25871_ (.A(_02604_),
    .B(_02616_),
    .S(_02588_),
    .Z(_02626_));
 MUX2_X1 _25872_ (.A(_02602_),
    .B(_02626_),
    .S(_02598_),
    .Z(_02627_));
 NAND2_X1 _25873_ (.A1(_02608_),
    .A2(_02620_),
    .ZN(_02628_));
 OAI22_X2 _25874_ (.A1(_02608_),
    .A2(_02625_),
    .B1(_02627_),
    .B2(_02628_),
    .ZN(_02629_));
 NAND2_X2 _25875_ (.A1(_02572_),
    .A2(_02629_),
    .ZN(_14124_));
 INV_X1 _25876_ (.A(_14124_),
    .ZN(_14119_));
 NAND2_X2 _25877_ (.A1(_02572_),
    .A2(_02620_),
    .ZN(_02630_));
 NOR2_X1 _25878_ (.A1(_02608_),
    .A2(_02630_),
    .ZN(_02631_));
 NAND2_X1 _25879_ (.A1(_02624_),
    .A2(_02631_),
    .ZN(_21763_));
 INV_X1 _25880_ (.A(_21763_),
    .ZN(_21767_));
 OR3_X1 _25881_ (.A1(_02608_),
    .A2(_02618_),
    .A3(_02630_),
    .ZN(_21756_));
 INV_X1 _25882_ (.A(_21756_),
    .ZN(_21760_));
 NOR2_X1 _25883_ (.A1(_02597_),
    .A2(_02587_),
    .ZN(_02632_));
 AND2_X1 _25884_ (.A1(_02597_),
    .A2(_02587_),
    .ZN(_02633_));
 AOI22_X2 _25885_ (.A1(_02616_),
    .A2(_02632_),
    .B1(_02633_),
    .B2(_02614_),
    .ZN(_02634_));
 NOR2_X4 _25886_ (.A1(_02598_),
    .A2(_02587_),
    .ZN(_02635_));
 NAND2_X1 _25887_ (.A1(_02601_),
    .A2(_02635_),
    .ZN(_02636_));
 AND2_X1 _25888_ (.A1(_02634_),
    .A2(_02636_),
    .ZN(_02637_));
 NAND2_X1 _25889_ (.A1(_02631_),
    .A2(_02637_),
    .ZN(_21791_));
 INV_X1 _25890_ (.A(_21791_),
    .ZN(_21795_));
 OR2_X1 _25891_ (.A1(_02598_),
    .A2(_02587_),
    .ZN(_02638_));
 MUX2_X1 _25892_ (.A(_02601_),
    .B(_02604_),
    .S(_02597_),
    .Z(_02639_));
 NOR2_X1 _25893_ (.A1(_02588_),
    .A2(_02639_),
    .ZN(_02640_));
 AOI21_X1 _25894_ (.A(_02640_),
    .B1(_02617_),
    .B2(_02588_),
    .ZN(_02641_));
 MUX2_X1 _25895_ (.A(_02638_),
    .B(_02641_),
    .S(_02611_),
    .Z(_02642_));
 OR2_X1 _25896_ (.A1(_02630_),
    .A2(_02642_),
    .ZN(_21770_));
 INV_X1 _25897_ (.A(_21770_),
    .ZN(_21774_));
 NOR2_X1 _25898_ (.A1(_02608_),
    .A2(_02627_),
    .ZN(_02643_));
 AOI21_X1 _25899_ (.A(_02643_),
    .B1(_02624_),
    .B2(_02608_),
    .ZN(_02644_));
 NOR2_X1 _25900_ (.A1(_02630_),
    .A2(_02644_),
    .ZN(_21777_));
 INV_X1 _25901_ (.A(_21777_),
    .ZN(_21781_));
 MUX2_X1 _25902_ (.A(_02618_),
    .B(_02606_),
    .S(_02611_),
    .Z(_02645_));
 NOR2_X1 _25903_ (.A1(_02630_),
    .A2(_02645_),
    .ZN(_21784_));
 INV_X1 _25904_ (.A(_21784_),
    .ZN(_21788_));
 NAND2_X1 _25905_ (.A1(_02634_),
    .A2(_02636_),
    .ZN(_02646_));
 MUX2_X1 _25906_ (.A(_00539_),
    .B(_00541_),
    .S(_02587_),
    .Z(_02647_));
 MUX2_X1 _25907_ (.A(_00535_),
    .B(_00538_),
    .S(_02587_),
    .Z(_02648_));
 MUX2_X1 _25908_ (.A(_02647_),
    .B(_02648_),
    .S(_02597_),
    .Z(_02649_));
 MUX2_X1 _25909_ (.A(_21724_),
    .B(_21718_),
    .S(_02587_),
    .Z(_02650_));
 MUX2_X1 _25910_ (.A(_21727_),
    .B(_21721_),
    .S(_02587_),
    .Z(_02651_));
 MUX2_X1 _25911_ (.A(_02650_),
    .B(_02651_),
    .S(_02597_),
    .Z(_02652_));
 MUX2_X1 _25912_ (.A(_02649_),
    .B(_02652_),
    .S(_02532_),
    .Z(_02653_));
 MUX2_X1 _25913_ (.A(_02646_),
    .B(_02653_),
    .S(_02611_),
    .Z(_02654_));
 NOR2_X1 _25914_ (.A1(_02630_),
    .A2(_02654_),
    .ZN(_21801_));
 INV_X1 _25915_ (.A(_21801_),
    .ZN(_21805_));
 NAND3_X1 _25916_ (.A1(_02611_),
    .A2(_02584_),
    .A3(_02635_),
    .ZN(_02655_));
 MUX2_X1 _25917_ (.A(_02591_),
    .B(_02600_),
    .S(_02588_),
    .Z(_02656_));
 MUX2_X1 _25918_ (.A(_02621_),
    .B(_02656_),
    .S(_02598_),
    .Z(_02657_));
 MUX2_X1 _25919_ (.A(_02641_),
    .B(_02657_),
    .S(_02611_),
    .Z(_02658_));
 OAI21_X1 _25920_ (.A(_02655_),
    .B1(_02658_),
    .B2(_02584_),
    .ZN(_02659_));
 NAND2_X1 _25921_ (.A1(_02572_),
    .A2(_02659_),
    .ZN(_21798_));
 INV_X1 _25922_ (.A(_21798_),
    .ZN(_21752_));
 XOR2_X2 _25923_ (.A(\g_reduce0[6].adder.b[15] ),
    .B(\g_reduce0[6].adder.a[15] ),
    .Z(_02660_));
 BUF_X4 _25924_ (.A(_02660_),
    .Z(_02661_));
 BUF_X2 _25925_ (.A(_21766_),
    .Z(_02662_));
 INV_X2 _25926_ (.A(_02662_),
    .ZN(_02663_));
 BUF_X2 _25927_ (.A(_21759_),
    .Z(_02664_));
 BUF_X4 _25928_ (.A(_21773_),
    .Z(_02665_));
 CLKBUF_X2 _25929_ (.A(_21780_),
    .Z(_02666_));
 NOR2_X1 _25930_ (.A1(_02666_),
    .A2(_21779_),
    .ZN(_02667_));
 NOR3_X1 _25931_ (.A1(_02665_),
    .A2(_21794_),
    .A3(_02667_),
    .ZN(_02668_));
 INV_X1 _25932_ (.A(_21786_),
    .ZN(_02669_));
 AOI21_X2 _25933_ (.A(_21748_),
    .B1(_14118_),
    .B2(_21749_),
    .ZN(_02670_));
 BUF_X2 _25934_ (.A(_21787_),
    .Z(_02671_));
 BUF_X4 _25935_ (.A(_21804_),
    .Z(_02672_));
 BUF_X1 _25936_ (.A(_21755_),
    .Z(_02673_));
 NAND3_X1 _25937_ (.A1(_02671_),
    .A2(_02672_),
    .A3(_02673_),
    .ZN(_02674_));
 AOI21_X1 _25938_ (.A(_21803_),
    .B1(_02672_),
    .B2(_21754_),
    .ZN(_02675_));
 INV_X2 _25939_ (.A(_02671_),
    .ZN(_02676_));
 OAI221_X1 _25940_ (.A(_02669_),
    .B1(_02670_),
    .B2(_02674_),
    .C1(_02675_),
    .C2(_02676_),
    .ZN(_02677_));
 OAI21_X1 _25941_ (.A(_02668_),
    .B1(_02677_),
    .B2(_21779_),
    .ZN(_02678_));
 INV_X2 _25942_ (.A(_21794_),
    .ZN(_02679_));
 AOI21_X1 _25943_ (.A(_21796_),
    .B1(_21775_),
    .B2(_02679_),
    .ZN(_02680_));
 AOI21_X1 _25944_ (.A(_02664_),
    .B1(_02678_),
    .B2(_02680_),
    .ZN(_02681_));
 OAI21_X2 _25945_ (.A(_02663_),
    .B1(_02681_),
    .B2(_21761_),
    .ZN(_02682_));
 INV_X1 _25946_ (.A(_21768_),
    .ZN(_02683_));
 AOI21_X4 _25947_ (.A(_02661_),
    .B1(_02682_),
    .B2(_02683_),
    .ZN(_02684_));
 OR4_X2 _25948_ (.A1(_02500_),
    .A2(_02607_),
    .A3(_02583_),
    .A4(_02638_),
    .ZN(_02685_));
 AND3_X1 _25949_ (.A1(_02495_),
    .A2(_02567_),
    .A3(_02570_),
    .ZN(_02686_));
 NAND4_X2 _25950_ (.A1(_02611_),
    .A2(_02583_),
    .A3(_02686_),
    .A4(_02635_),
    .ZN(_02687_));
 OAI211_X2 _25951_ (.A(_02493_),
    .B(_02547_),
    .C1(_02560_),
    .C2(_02499_),
    .ZN(_02688_));
 MUX2_X1 _25952_ (.A(_02688_),
    .B(_02493_),
    .S(_02583_),
    .Z(_02689_));
 NAND3_X2 _25953_ (.A1(_02552_),
    .A2(_02611_),
    .A3(_02635_),
    .ZN(_02690_));
 OAI211_X4 _25954_ (.A(_02685_),
    .B(_02687_),
    .C1(_02689_),
    .C2(_02690_),
    .ZN(_02691_));
 BUF_X2 _25955_ (.A(_21758_),
    .Z(_02692_));
 INV_X1 _25956_ (.A(_02692_),
    .ZN(_02693_));
 BUF_X2 _25957_ (.A(_21793_),
    .Z(_02694_));
 OR2_X2 _25958_ (.A1(_21782_),
    .A2(_21789_),
    .ZN(_02695_));
 OR3_X1 _25959_ (.A1(_21772_),
    .A2(_02676_),
    .A3(_02695_),
    .ZN(_02696_));
 INV_X1 _25960_ (.A(_02665_),
    .ZN(_02697_));
 INV_X1 _25961_ (.A(_21782_),
    .ZN(_02698_));
 AOI21_X2 _25962_ (.A(_02697_),
    .B1(_02698_),
    .B2(_02666_),
    .ZN(_02699_));
 OAI21_X2 _25963_ (.A(_02696_),
    .B1(_02699_),
    .B2(_21772_),
    .ZN(_02700_));
 NAND2_X1 _25964_ (.A1(_14123_),
    .A2(_21751_),
    .ZN(_02701_));
 NOR2_X1 _25965_ (.A1(_21750_),
    .A2(_21799_),
    .ZN(_02702_));
 INV_X1 _25966_ (.A(_21800_),
    .ZN(_02703_));
 INV_X1 _25967_ (.A(_21799_),
    .ZN(_02704_));
 AOI221_X2 _25968_ (.A(_02672_),
    .B1(_02701_),
    .B2(_02702_),
    .C1(_02703_),
    .C2(_02704_),
    .ZN(_02705_));
 NOR4_X4 _25969_ (.A1(_21772_),
    .A2(_21806_),
    .A3(_02705_),
    .A4(_02695_),
    .ZN(_02706_));
 NOR3_X4 _25970_ (.A1(_02679_),
    .A2(_02700_),
    .A3(_02706_),
    .ZN(_02707_));
 OAI21_X1 _25971_ (.A(_02664_),
    .B1(_02694_),
    .B2(_02707_),
    .ZN(_02708_));
 AOI21_X2 _25972_ (.A(_02663_),
    .B1(_02693_),
    .B2(_02708_),
    .ZN(_02709_));
 OAI21_X4 _25973_ (.A(_02661_),
    .B1(_02709_),
    .B2(_21765_),
    .ZN(_02710_));
 AOI21_X4 _25974_ (.A(_02684_),
    .B1(_02691_),
    .B2(_02710_),
    .ZN(_02711_));
 XNOR2_X2 _25975_ (.A(\g_reduce0[6].adder.b[15] ),
    .B(\g_reduce0[6].adder.a[15] ),
    .ZN(_02712_));
 BUF_X4 _25976_ (.A(_02712_),
    .Z(_02713_));
 BUF_X4 _25977_ (.A(_02713_),
    .Z(_02714_));
 NOR4_X4 _25978_ (.A1(_02694_),
    .A2(_02692_),
    .A3(_02714_),
    .A4(_02707_),
    .ZN(_02715_));
 AND2_X1 _25979_ (.A1(_02712_),
    .A2(_02680_),
    .ZN(_02716_));
 AOI221_X1 _25980_ (.A(_02664_),
    .B1(_02692_),
    .B2(_02660_),
    .C1(_02678_),
    .C2(_02716_),
    .ZN(_02717_));
 NAND2_X1 _25981_ (.A1(_21761_),
    .A2(_02713_),
    .ZN(_02718_));
 INV_X1 _25982_ (.A(_02718_),
    .ZN(_02719_));
 OR2_X1 _25983_ (.A1(_02717_),
    .A2(_02719_),
    .ZN(_02720_));
 OAI21_X1 _25984_ (.A(_02662_),
    .B1(_02715_),
    .B2(_02720_),
    .ZN(_02721_));
 OR4_X2 _25985_ (.A1(_02694_),
    .A2(_02692_),
    .A3(_02714_),
    .A4(_02707_),
    .ZN(_02722_));
 NOR2_X2 _25986_ (.A1(_02717_),
    .A2(_02719_),
    .ZN(_02723_));
 NAND3_X1 _25987_ (.A1(_02663_),
    .A2(_02722_),
    .A3(_02723_),
    .ZN(_02724_));
 INV_X1 _25988_ (.A(_21775_),
    .ZN(_02725_));
 AOI21_X1 _25989_ (.A(_21794_),
    .B1(_02725_),
    .B2(_02665_),
    .ZN(_02726_));
 OR2_X1 _25990_ (.A1(_21796_),
    .A2(_21775_),
    .ZN(_02727_));
 INV_X1 _25991_ (.A(_21779_),
    .ZN(_02728_));
 AOI21_X2 _25992_ (.A(_21754_),
    .B1(_14121_),
    .B2(_02673_),
    .ZN(_02729_));
 NAND3_X1 _25993_ (.A1(_02666_),
    .A2(_02671_),
    .A3(_02672_),
    .ZN(_02730_));
 AOI21_X1 _25994_ (.A(_21786_),
    .B1(_21803_),
    .B2(_02671_),
    .ZN(_02731_));
 INV_X1 _25995_ (.A(_02666_),
    .ZN(_02732_));
 OAI221_X2 _25996_ (.A(_02728_),
    .B1(_02729_),
    .B2(_02730_),
    .C1(_02731_),
    .C2(_02732_),
    .ZN(_02733_));
 OAI22_X2 _25997_ (.A1(_21796_),
    .A2(_02726_),
    .B1(_02727_),
    .B2(_02733_),
    .ZN(_02734_));
 OR3_X1 _25998_ (.A1(_02664_),
    .A2(_02660_),
    .A3(_02734_),
    .ZN(_02735_));
 NAND3_X1 _25999_ (.A1(_02664_),
    .A2(_02714_),
    .A3(_02734_),
    .ZN(_02736_));
 INV_X1 _26000_ (.A(_02664_),
    .ZN(_02737_));
 OR2_X1 _26001_ (.A1(_02694_),
    .A2(_21772_),
    .ZN(_02738_));
 OAI22_X2 _26002_ (.A1(_21794_),
    .A2(_02694_),
    .B1(_02699_),
    .B2(_02738_),
    .ZN(_02739_));
 INV_X1 _26003_ (.A(_21806_),
    .ZN(_02740_));
 AOI21_X1 _26004_ (.A(_21799_),
    .B1(_14125_),
    .B2(_21800_),
    .ZN(_02741_));
 OAI21_X2 _26005_ (.A(_02740_),
    .B1(_02741_),
    .B2(_02672_),
    .ZN(_02742_));
 AOI211_X2 _26006_ (.A(_02695_),
    .B(_02738_),
    .C1(_02742_),
    .C2(_02676_),
    .ZN(_02743_));
 OR4_X1 _26007_ (.A1(_02737_),
    .A2(_02713_),
    .A3(_02739_),
    .A4(_02743_),
    .ZN(_02744_));
 NOR2_X1 _26008_ (.A1(_02664_),
    .A2(_02713_),
    .ZN(_02745_));
 OAI21_X2 _26009_ (.A(_02745_),
    .B1(_02743_),
    .B2(_02739_),
    .ZN(_02746_));
 NAND4_X4 _26010_ (.A1(_02735_),
    .A2(_02736_),
    .A3(_02744_),
    .A4(_02746_),
    .ZN(_02747_));
 INV_X1 _26011_ (.A(_02747_),
    .ZN(_02748_));
 NAND3_X1 _26012_ (.A1(_02721_),
    .A2(_02724_),
    .A3(_02748_),
    .ZN(_02749_));
 NAND2_X1 _26013_ (.A1(_21765_),
    .A2(_02661_),
    .ZN(_02750_));
 NOR2_X1 _26014_ (.A1(_02663_),
    .A2(_02714_),
    .ZN(_02751_));
 NOR3_X1 _26015_ (.A1(_02737_),
    .A2(_02739_),
    .A3(_02743_),
    .ZN(_02752_));
 OAI21_X1 _26016_ (.A(_02751_),
    .B1(_02752_),
    .B2(_02692_),
    .ZN(_02753_));
 NOR3_X1 _26017_ (.A1(_02664_),
    .A2(_02662_),
    .A3(_02734_),
    .ZN(_02754_));
 INV_X1 _26018_ (.A(_21761_),
    .ZN(_02755_));
 OAI21_X1 _26019_ (.A(_02683_),
    .B1(_02755_),
    .B2(_02662_),
    .ZN(_02756_));
 OR3_X1 _26020_ (.A1(_02661_),
    .A2(_02754_),
    .A3(_02756_),
    .ZN(_02757_));
 AND3_X2 _26021_ (.A1(_02750_),
    .A2(_02753_),
    .A3(_02757_),
    .ZN(_02758_));
 AND2_X1 _26022_ (.A1(_02749_),
    .A2(_02758_),
    .ZN(_02759_));
 NAND3_X1 _26023_ (.A1(_02750_),
    .A2(_02753_),
    .A3(_02757_),
    .ZN(_02760_));
 AND2_X1 _26024_ (.A1(_02749_),
    .A2(_02760_),
    .ZN(_02761_));
 MUX2_X2 _26025_ (.A(_02759_),
    .B(_02761_),
    .S(_02691_),
    .Z(_02762_));
 AOI21_X4 _26026_ (.A(_02663_),
    .B1(_02722_),
    .B2(_02723_),
    .ZN(_02763_));
 NOR3_X4 _26027_ (.A1(_02662_),
    .A2(_02715_),
    .A3(_02720_),
    .ZN(_02764_));
 NOR2_X1 _26028_ (.A1(_02763_),
    .A2(_02764_),
    .ZN(_02765_));
 OR3_X2 _26029_ (.A1(_02713_),
    .A2(_02700_),
    .A3(_02706_),
    .ZN(_02766_));
 NOR2_X1 _26030_ (.A1(_02665_),
    .A2(_02667_),
    .ZN(_02767_));
 OAI21_X1 _26031_ (.A(_02767_),
    .B1(_02677_),
    .B2(_21779_),
    .ZN(_02768_));
 NAND3_X2 _26032_ (.A1(_02725_),
    .A2(_02714_),
    .A3(_02768_),
    .ZN(_02769_));
 AND3_X2 _26033_ (.A1(_02679_),
    .A2(_02766_),
    .A3(_02769_),
    .ZN(_02770_));
 AOI21_X4 _26034_ (.A(_02679_),
    .B1(_02766_),
    .B2(_02769_),
    .ZN(_02771_));
 OAI21_X2 _26035_ (.A(_02676_),
    .B1(_21806_),
    .B2(_02705_),
    .ZN(_02772_));
 NOR2_X1 _26036_ (.A1(_21789_),
    .A2(_02713_),
    .ZN(_02773_));
 AOI22_X4 _26037_ (.A1(_02713_),
    .A2(_02677_),
    .B1(_02772_),
    .B2(_02773_),
    .ZN(_02774_));
 XNOR2_X2 _26038_ (.A(_02666_),
    .B(_02774_),
    .ZN(_02775_));
 INV_X1 _26039_ (.A(_02672_),
    .ZN(_02776_));
 INV_X1 _26040_ (.A(_02673_),
    .ZN(_02777_));
 NOR2_X1 _26041_ (.A1(_02777_),
    .A2(_02670_),
    .ZN(_02778_));
 OAI21_X1 _26042_ (.A(_02712_),
    .B1(_02778_),
    .B2(_21754_),
    .ZN(_02779_));
 AOI21_X1 _26043_ (.A(_21750_),
    .B1(_14123_),
    .B2(_21751_),
    .ZN(_02780_));
 OAI21_X1 _26044_ (.A(_02704_),
    .B1(_02703_),
    .B2(_02780_),
    .ZN(_02781_));
 OAI21_X1 _26045_ (.A(_02779_),
    .B1(_02781_),
    .B2(_02713_),
    .ZN(_02782_));
 XNOR2_X2 _26046_ (.A(_02776_),
    .B(_02782_),
    .ZN(_02783_));
 NOR2_X1 _26047_ (.A1(_02676_),
    .A2(_02660_),
    .ZN(_02784_));
 NOR2_X1 _26048_ (.A1(_02671_),
    .A2(_02660_),
    .ZN(_02785_));
 INV_X1 _26049_ (.A(_21803_),
    .ZN(_02786_));
 OAI21_X1 _26050_ (.A(_02786_),
    .B1(_02729_),
    .B2(_02776_),
    .ZN(_02787_));
 MUX2_X1 _26051_ (.A(_02784_),
    .B(_02785_),
    .S(_02787_),
    .Z(_02788_));
 NOR2_X1 _26052_ (.A1(_02671_),
    .A2(_02713_),
    .ZN(_02789_));
 NOR2_X1 _26053_ (.A1(_02676_),
    .A2(_02713_),
    .ZN(_02790_));
 MUX2_X1 _26054_ (.A(_02789_),
    .B(_02790_),
    .S(_02742_),
    .Z(_02791_));
 NOR2_X2 _26055_ (.A1(_02788_),
    .A2(_02791_),
    .ZN(_02792_));
 AOI21_X1 _26056_ (.A(_02775_),
    .B1(_02783_),
    .B2(_02792_),
    .ZN(_02793_));
 NAND2_X1 _26057_ (.A1(_21782_),
    .A2(_02660_),
    .ZN(_02794_));
 NAND2_X1 _26058_ (.A1(_02732_),
    .A2(_02660_),
    .ZN(_02795_));
 AOI21_X1 _26059_ (.A(_21789_),
    .B1(_02742_),
    .B2(_02676_),
    .ZN(_02796_));
 OAI221_X2 _26060_ (.A(_02794_),
    .B1(_02795_),
    .B2(_02796_),
    .C1(_02660_),
    .C2(_02733_),
    .ZN(_02797_));
 XNOR2_X2 _26061_ (.A(_02697_),
    .B(_02797_),
    .ZN(_02798_));
 OAI221_X1 _26062_ (.A(_02765_),
    .B1(_02770_),
    .B2(_02771_),
    .C1(_02793_),
    .C2(_02798_),
    .ZN(_02799_));
 BUF_X1 _26063_ (.A(_02799_),
    .Z(_02800_));
 XNOR2_X1 _26064_ (.A(_14121_),
    .B(_02673_),
    .ZN(_02801_));
 XNOR2_X1 _26065_ (.A(_14125_),
    .B(_21800_),
    .ZN(_02802_));
 MUX2_X1 _26066_ (.A(_02801_),
    .B(_02802_),
    .S(_02660_),
    .Z(_02803_));
 CLKBUF_X3 _26067_ (.A(_02803_),
    .Z(_02804_));
 NAND2_X2 _26068_ (.A1(_02792_),
    .A2(_02804_),
    .ZN(_02805_));
 OR2_X1 _26069_ (.A1(_02798_),
    .A2(_02805_),
    .ZN(_02806_));
 NOR2_X1 _26070_ (.A1(_21810_),
    .A2(_02661_),
    .ZN(_02807_));
 INV_X1 _26071_ (.A(_02807_),
    .ZN(_02808_));
 NOR4_X1 _26072_ (.A1(_02611_),
    .A2(_02653_),
    .A3(_02806_),
    .A4(_02808_),
    .ZN(_02809_));
 AND3_X2 _26073_ (.A1(_02561_),
    .A2(_02566_),
    .A3(_02571_),
    .ZN(_02810_));
 NOR2_X1 _26074_ (.A1(_02810_),
    .A2(_02584_),
    .ZN(_02811_));
 AOI21_X1 _26075_ (.A(_02800_),
    .B1(_02809_),
    .B2(_02811_),
    .ZN(_02812_));
 OR3_X1 _26076_ (.A1(_21812_),
    .A2(_02714_),
    .A3(_02806_),
    .ZN(_02813_));
 NAND3_X1 _26077_ (.A1(_02610_),
    .A2(_02634_),
    .A3(_02636_),
    .ZN(_02814_));
 NOR3_X1 _26078_ (.A1(_02506_),
    .A2(_21736_),
    .A3(_21744_),
    .ZN(_02815_));
 NOR3_X1 _26079_ (.A1(_02597_),
    .A2(_00533_),
    .A3(_21744_),
    .ZN(_02816_));
 MUX2_X1 _26080_ (.A(_02815_),
    .B(_02816_),
    .S(_02531_),
    .Z(_02817_));
 INV_X1 _26081_ (.A(_02613_),
    .ZN(_02818_));
 INV_X1 _26082_ (.A(_00536_),
    .ZN(_02819_));
 INV_X1 _26083_ (.A(_21730_),
    .ZN(_02820_));
 MUX2_X1 _26084_ (.A(_02819_),
    .B(_02820_),
    .S(_02532_),
    .Z(_02821_));
 AOI221_X2 _26085_ (.A(_02817_),
    .B1(_02633_),
    .B2(_02595_),
    .C1(_02818_),
    .C2(_02821_),
    .ZN(_02822_));
 MUX2_X1 _26086_ (.A(_02653_),
    .B(_02822_),
    .S(_02610_),
    .Z(_02823_));
 MUX2_X1 _26087_ (.A(_02814_),
    .B(_02823_),
    .S(_02620_),
    .Z(_02824_));
 NOR2_X1 _26088_ (.A1(_02810_),
    .A2(_02824_),
    .ZN(_02825_));
 AND2_X1 _26089_ (.A1(_14122_),
    .A2(_02714_),
    .ZN(_02826_));
 AOI21_X2 _26090_ (.A(_02826_),
    .B1(_02661_),
    .B2(_14126_),
    .ZN(_02827_));
 AOI21_X1 _26091_ (.A(_02817_),
    .B1(_02821_),
    .B2(_02818_),
    .ZN(_02828_));
 NAND2_X1 _26092_ (.A1(_02595_),
    .A2(_02633_),
    .ZN(_02829_));
 NAND2_X1 _26093_ (.A1(_02828_),
    .A2(_02829_),
    .ZN(_02830_));
 MUX2_X1 _26094_ (.A(_02637_),
    .B(_02830_),
    .S(_02620_),
    .Z(_02831_));
 NOR3_X1 _26095_ (.A1(_02810_),
    .A2(_02608_),
    .A3(_02808_),
    .ZN(_02832_));
 AOI21_X1 _26096_ (.A(_02827_),
    .B1(_02831_),
    .B2(_02832_),
    .ZN(_02833_));
 OAI221_X2 _26097_ (.A(_02812_),
    .B1(_02813_),
    .B2(_02825_),
    .C1(_02806_),
    .C2(_02833_),
    .ZN(_02834_));
 BUF_X4 _26098_ (.A(_02834_),
    .Z(_02835_));
 NAND2_X2 _26099_ (.A1(_02762_),
    .A2(_02835_),
    .ZN(_02836_));
 NAND2_X2 _26100_ (.A1(_02711_),
    .A2(_02836_),
    .ZN(_21814_));
 INV_X2 _26101_ (.A(_21814_),
    .ZN(_21816_));
 NOR3_X4 _26102_ (.A1(_02805_),
    .A2(_02775_),
    .A3(_02783_),
    .ZN(_02837_));
 XNOR2_X2 _26103_ (.A(_02665_),
    .B(_02797_),
    .ZN(_02838_));
 OAI211_X4 _26104_ (.A(_02747_),
    .B(_02838_),
    .C1(_02770_),
    .C2(_02771_),
    .ZN(_02839_));
 NOR4_X4 _26105_ (.A1(_02763_),
    .A2(_02764_),
    .A3(_02837_),
    .A4(_02839_),
    .ZN(_02840_));
 NOR3_X1 _26106_ (.A1(_02710_),
    .A2(_02758_),
    .A3(_02840_),
    .ZN(_02841_));
 OR2_X1 _26107_ (.A1(_02684_),
    .A2(_02760_),
    .ZN(_02842_));
 NOR2_X1 _26108_ (.A1(_02840_),
    .A2(_02842_),
    .ZN(_02843_));
 NOR4_X1 _26109_ (.A1(_02500_),
    .A2(_02608_),
    .A3(_02583_),
    .A4(_02638_),
    .ZN(_02844_));
 AND4_X1 _26110_ (.A1(_02610_),
    .A2(_02583_),
    .A3(_02686_),
    .A4(_02635_),
    .ZN(_02845_));
 AOI211_X2 _26111_ (.A(_02567_),
    .B(_02565_),
    .C1(_02562_),
    .C2(_02498_),
    .ZN(_02846_));
 MUX2_X1 _26112_ (.A(_02846_),
    .B(_02567_),
    .S(_02583_),
    .Z(_02847_));
 AND3_X1 _26113_ (.A1(_02552_),
    .A2(_02610_),
    .A3(_02635_),
    .ZN(_02848_));
 AOI211_X2 _26114_ (.A(_02844_),
    .B(_02845_),
    .C1(_02847_),
    .C2(_02848_),
    .ZN(_02849_));
 MUX2_X1 _26115_ (.A(_02841_),
    .B(_02843_),
    .S(_02849_),
    .Z(_02850_));
 XNOR2_X2 _26116_ (.A(_21819_),
    .B(_02850_),
    .ZN(_02851_));
 INV_X4 _26117_ (.A(_02851_),
    .ZN(_02852_));
 BUF_X8 _26118_ (.A(_02852_),
    .Z(_21840_));
 OR2_X1 _26119_ (.A1(_02710_),
    .A2(_02758_),
    .ZN(_02853_));
 MUX2_X1 _26120_ (.A(_02842_),
    .B(_02853_),
    .S(_02691_),
    .Z(_02854_));
 BUF_X4 _26121_ (.A(_02854_),
    .Z(_02855_));
 CLKBUF_X3 _26122_ (.A(_21815_),
    .Z(_02856_));
 MUX2_X2 _26123_ (.A(_21810_),
    .B(_21812_),
    .S(_02661_),
    .Z(_02857_));
 NAND2_X1 _26124_ (.A1(_02856_),
    .A2(_02857_),
    .ZN(_02858_));
 OAI21_X1 _26125_ (.A(_02714_),
    .B1(_02824_),
    .B2(_02810_),
    .ZN(_02859_));
 NOR3_X1 _26126_ (.A1(_02810_),
    .A2(_02584_),
    .A3(_02823_),
    .ZN(_02860_));
 NOR3_X1 _26127_ (.A1(_02810_),
    .A2(_02620_),
    .A3(_02814_),
    .ZN(_02861_));
 OAI21_X1 _26128_ (.A(_02661_),
    .B1(_02860_),
    .B2(_02861_),
    .ZN(_02862_));
 NAND2_X1 _26129_ (.A1(_02859_),
    .A2(_02862_),
    .ZN(_02863_));
 OAI21_X1 _26130_ (.A(_02858_),
    .B1(_02863_),
    .B2(_02856_),
    .ZN(_02864_));
 NAND2_X1 _26131_ (.A1(_02855_),
    .A2(_02864_),
    .ZN(_02865_));
 NAND2_X2 _26132_ (.A1(_02721_),
    .A2(_02724_),
    .ZN(_02866_));
 OR2_X2 _26133_ (.A1(_02866_),
    .A2(_02839_),
    .ZN(_02867_));
 OR2_X2 _26134_ (.A1(_02788_),
    .A2(_02791_),
    .ZN(_02868_));
 XNOR2_X2 _26135_ (.A(_02732_),
    .B(_02774_),
    .ZN(_02869_));
 OAI21_X1 _26136_ (.A(_02804_),
    .B1(_02827_),
    .B2(_02857_),
    .ZN(_02870_));
 OAI21_X1 _26137_ (.A(_02869_),
    .B1(_02783_),
    .B2(_02870_),
    .ZN(_02871_));
 OR2_X1 _26138_ (.A1(_02868_),
    .A2(_02871_),
    .ZN(_02872_));
 NOR2_X2 _26139_ (.A1(_02867_),
    .A2(_02872_),
    .ZN(_02873_));
 NOR2_X2 _26140_ (.A1(_02867_),
    .A2(_02840_),
    .ZN(_02874_));
 OR3_X2 _26141_ (.A1(_02854_),
    .A2(_02873_),
    .A3(_02874_),
    .ZN(_02875_));
 BUF_X4 _26142_ (.A(_02762_),
    .Z(_02876_));
 NOR2_X1 _26143_ (.A1(_02684_),
    .A2(_02760_),
    .ZN(_02877_));
 NOR2_X1 _26144_ (.A1(_02710_),
    .A2(_02758_),
    .ZN(_02878_));
 MUX2_X2 _26145_ (.A(_02877_),
    .B(_02878_),
    .S(_02691_),
    .Z(_02879_));
 NAND3_X2 _26146_ (.A1(_02876_),
    .A2(_02800_),
    .A3(_02879_),
    .ZN(_02880_));
 AOI21_X4 _26147_ (.A(_02851_),
    .B1(_02875_),
    .B2(_02880_),
    .ZN(_02881_));
 BUF_X1 _26148_ (.A(_14128_),
    .Z(_02882_));
 NAND2_X2 _26149_ (.A1(_02882_),
    .A2(_02711_),
    .ZN(_02883_));
 AOI22_X2 _26150_ (.A1(_02762_),
    .A2(_02800_),
    .B1(_02859_),
    .B2(_02862_),
    .ZN(_02884_));
 NOR2_X1 _26151_ (.A1(_02798_),
    .A2(_02805_),
    .ZN(_02885_));
 MUX2_X2 _26152_ (.A(_14126_),
    .B(_14122_),
    .S(_02714_),
    .Z(_02886_));
 NOR2_X1 _26153_ (.A1(_02653_),
    .A2(_02808_),
    .ZN(_02887_));
 NAND4_X2 _26154_ (.A1(_02572_),
    .A2(_02608_),
    .A3(_02620_),
    .A4(_02887_),
    .ZN(_02888_));
 NAND3_X1 _26155_ (.A1(_02572_),
    .A2(_02611_),
    .A3(_02807_),
    .ZN(_02889_));
 MUX2_X1 _26156_ (.A(_02646_),
    .B(_02822_),
    .S(_02620_),
    .Z(_02890_));
 OAI211_X2 _26157_ (.A(_02886_),
    .B(_02888_),
    .C1(_02889_),
    .C2(_02890_),
    .ZN(_02891_));
 NAND3_X1 _26158_ (.A1(_02762_),
    .A2(_02885_),
    .A3(_02891_),
    .ZN(_02892_));
 AOI21_X2 _26159_ (.A(_02883_),
    .B1(_02884_),
    .B2(_02892_),
    .ZN(_02893_));
 NAND2_X1 _26160_ (.A1(_02881_),
    .A2(_02893_),
    .ZN(_02894_));
 NAND2_X1 _26161_ (.A1(_02856_),
    .A2(_02886_),
    .ZN(_02895_));
 XNOR2_X2 _26162_ (.A(_02691_),
    .B(_02758_),
    .ZN(_02896_));
 AND2_X1 _26163_ (.A1(_02683_),
    .A2(_02682_),
    .ZN(_02897_));
 INV_X1 _26164_ (.A(_02710_),
    .ZN(_02898_));
 OAI22_X4 _26165_ (.A1(_02661_),
    .A2(_02897_),
    .B1(_02849_),
    .B2(_02898_),
    .ZN(_02899_));
 OAI221_X2 _26166_ (.A(_02895_),
    .B1(_02896_),
    .B2(_02899_),
    .C1(_02856_),
    .C2(_02857_),
    .ZN(_02900_));
 AND2_X1 _26167_ (.A1(_21810_),
    .A2(_02714_),
    .ZN(_02901_));
 AOI21_X2 _26168_ (.A(_02901_),
    .B1(_02661_),
    .B2(_21812_),
    .ZN(_02902_));
 CLKBUF_X3 _26169_ (.A(_02882_),
    .Z(_02903_));
 AOI22_X2 _26170_ (.A1(_02876_),
    .A2(_02835_),
    .B1(_02902_),
    .B2(_02903_),
    .ZN(_02904_));
 INV_X1 _26171_ (.A(_02882_),
    .ZN(_02905_));
 CLKBUF_X3 _26172_ (.A(_02905_),
    .Z(_02906_));
 XNOR2_X2 _26173_ (.A(_02849_),
    .B(_02758_),
    .ZN(_02907_));
 NAND2_X2 _26174_ (.A1(_02749_),
    .A2(_02907_),
    .ZN(_02908_));
 OAI33_X1 _26175_ (.A1(_02860_),
    .A2(_02861_),
    .A3(_02813_),
    .B1(_02888_),
    .B2(_02798_),
    .B3(_02805_),
    .ZN(_02909_));
 OAI21_X1 _26176_ (.A(_02886_),
    .B1(_02890_),
    .B2(_02889_),
    .ZN(_02910_));
 AOI211_X2 _26177_ (.A(_02800_),
    .B(_02909_),
    .C1(_02885_),
    .C2(_02910_),
    .ZN(_02911_));
 NOR4_X2 _26178_ (.A1(_02906_),
    .A2(_02908_),
    .A3(_02911_),
    .A4(_02863_),
    .ZN(_02912_));
 OAI21_X1 _26179_ (.A(_02881_),
    .B1(_02904_),
    .B2(_02912_),
    .ZN(_02913_));
 AOI22_X2 _26180_ (.A1(_02865_),
    .A2(_02894_),
    .B1(_02900_),
    .B2(_02913_),
    .ZN(_21821_));
 NOR4_X4 _26181_ (.A1(_02482_),
    .A2(_02483_),
    .A3(_02484_),
    .A4(_02485_),
    .ZN(_02914_));
 NAND2_X1 _26182_ (.A1(\g_reduce0[6].adder.b[0] ),
    .A2(_02914_),
    .ZN(_02915_));
 BUF_X4 _26183_ (.A(_02486_),
    .Z(_02916_));
 OR4_X1 _26184_ (.A1(_02487_),
    .A2(_02488_),
    .A3(_02489_),
    .A4(_02490_),
    .ZN(_02917_));
 BUF_X4 _26185_ (.A(_02917_),
    .Z(_02918_));
 OAI21_X1 _26186_ (.A(_02916_),
    .B1(_02918_),
    .B2(\g_reduce0[6].adder.a[0] ),
    .ZN(_02919_));
 BUF_X4 _26187_ (.A(_02856_),
    .Z(_02920_));
 BUF_X4 _26188_ (.A(_02879_),
    .Z(_02921_));
 NAND2_X1 _26189_ (.A1(_02921_),
    .A2(_02874_),
    .ZN(_02922_));
 NAND2_X2 _26190_ (.A1(_02921_),
    .A2(_02873_),
    .ZN(_02923_));
 OAI211_X4 _26191_ (.A(_02711_),
    .B(_02922_),
    .C1(_02923_),
    .C2(_02835_),
    .ZN(_02924_));
 INV_X2 _26192_ (.A(_02924_),
    .ZN(_21844_));
 NOR2_X1 _26193_ (.A1(_02882_),
    .A2(_02886_),
    .ZN(_02925_));
 AOI21_X1 _26194_ (.A(_02925_),
    .B1(_02783_),
    .B2(_02903_),
    .ZN(_02926_));
 NOR2_X1 _26195_ (.A1(_02899_),
    .A2(_02926_),
    .ZN(_02927_));
 NAND2_X1 _26196_ (.A1(_02836_),
    .A2(_02927_),
    .ZN(_02928_));
 NAND2_X1 _26197_ (.A1(_02906_),
    .A2(_02857_),
    .ZN(_02929_));
 OAI21_X1 _26198_ (.A(_02929_),
    .B1(_02804_),
    .B2(_02906_),
    .ZN(_02930_));
 NAND4_X1 _26199_ (.A1(_02711_),
    .A2(_02876_),
    .A3(_02835_),
    .A4(_02930_),
    .ZN(_02931_));
 AND2_X1 _26200_ (.A1(_02928_),
    .A2(_02931_),
    .ZN(_02932_));
 OAI221_X2 _26201_ (.A(_02711_),
    .B1(_02763_),
    .B2(_02764_),
    .C1(_02748_),
    .C2(_02896_),
    .ZN(_02933_));
 OAI221_X2 _26202_ (.A(_21840_),
    .B1(_21844_),
    .B2(_02932_),
    .C1(_02933_),
    .C2(_02903_),
    .ZN(_02934_));
 NOR2_X1 _26203_ (.A1(_02903_),
    .A2(_02899_),
    .ZN(_02935_));
 NAND4_X1 _26204_ (.A1(_02876_),
    .A2(_02868_),
    .A3(_02835_),
    .A4(_02935_),
    .ZN(_02936_));
 NOR2_X1 _26205_ (.A1(_02770_),
    .A2(_02771_),
    .ZN(_02937_));
 NOR2_X1 _26206_ (.A1(_02765_),
    .A2(_02896_),
    .ZN(_02938_));
 OAI221_X2 _26207_ (.A(_02711_),
    .B1(_02908_),
    .B2(_02798_),
    .C1(_02937_),
    .C2(_02938_),
    .ZN(_02939_));
 NOR2_X1 _26208_ (.A1(_02908_),
    .A2(_02911_),
    .ZN(_02940_));
 NAND2_X1 _26209_ (.A1(_02775_),
    .A2(_02935_),
    .ZN(_02941_));
 OAI221_X2 _26210_ (.A(_02936_),
    .B1(_02939_),
    .B2(_02906_),
    .C1(_02940_),
    .C2(_02941_),
    .ZN(_02942_));
 AND2_X1 _26211_ (.A1(_02893_),
    .A2(_02924_),
    .ZN(_02943_));
 OR2_X1 _26212_ (.A1(_02942_),
    .A2(_02943_),
    .ZN(_02944_));
 OAI21_X2 _26213_ (.A(_02934_),
    .B1(_02944_),
    .B2(_21840_),
    .ZN(_02945_));
 OAI22_X4 _26214_ (.A1(_02920_),
    .A2(_02711_),
    .B1(_02855_),
    .B2(_02945_),
    .ZN(_02946_));
 NAND2_X1 _26215_ (.A1(_02906_),
    .A2(_02711_),
    .ZN(_02947_));
 NOR2_X1 _26216_ (.A1(_02851_),
    .A2(_02947_),
    .ZN(_02948_));
 INV_X1 _26217_ (.A(_02863_),
    .ZN(_02949_));
 MUX2_X2 _26218_ (.A(_02949_),
    .B(_02857_),
    .S(_21816_),
    .Z(_02950_));
 OAI21_X1 _26219_ (.A(_02876_),
    .B1(_02885_),
    .B2(_02800_),
    .ZN(_02951_));
 AND2_X1 _26220_ (.A1(_02804_),
    .A2(_02951_),
    .ZN(_02952_));
 AND2_X1 _26221_ (.A1(_02762_),
    .A2(_02800_),
    .ZN(_02953_));
 OR3_X1 _26222_ (.A1(_02899_),
    .A2(_02804_),
    .A3(_02953_),
    .ZN(_02954_));
 AOI22_X4 _26223_ (.A1(_02711_),
    .A2(_02952_),
    .B1(_02954_),
    .B2(_02886_),
    .ZN(_02955_));
 NOR2_X1 _26224_ (.A1(_02851_),
    .A2(_02883_),
    .ZN(_02956_));
 AOI222_X2 _26225_ (.A1(_21817_),
    .A2(_02851_),
    .B1(_02948_),
    .B2(_02950_),
    .C1(_02955_),
    .C2(_02956_),
    .ZN(_02957_));
 NOR2_X1 _26226_ (.A1(_02856_),
    .A2(_02899_),
    .ZN(_02958_));
 INV_X1 _26227_ (.A(_02958_),
    .ZN(_02959_));
 NAND2_X1 _26228_ (.A1(_02856_),
    .A2(_02907_),
    .ZN(_02960_));
 AOI211_X4 _26229_ (.A(_21844_),
    .B(_02957_),
    .C1(_02959_),
    .C2(_02960_),
    .ZN(_02961_));
 NOR3_X1 _26230_ (.A1(_02866_),
    .A2(_02896_),
    .A3(_02851_),
    .ZN(_02962_));
 NOR2_X1 _26231_ (.A1(_02849_),
    .A2(_02898_),
    .ZN(_02963_));
 NOR4_X1 _26232_ (.A1(_02684_),
    .A2(_02963_),
    .A3(_02876_),
    .A4(_02838_),
    .ZN(_02964_));
 NOR2_X1 _26233_ (.A1(_02838_),
    .A2(_02800_),
    .ZN(_02965_));
 OAI33_X1 _26234_ (.A1(_02899_),
    .A2(_02876_),
    .A3(_02798_),
    .B1(_02775_),
    .B2(_02964_),
    .B3(_02965_),
    .ZN(_02966_));
 AOI21_X1 _26235_ (.A(_02962_),
    .B1(_02966_),
    .B2(_02851_),
    .ZN(_02967_));
 NOR2_X1 _26236_ (.A1(_02906_),
    .A2(_02967_),
    .ZN(_02968_));
 NAND2_X1 _26237_ (.A1(_21844_),
    .A2(_02958_),
    .ZN(_02969_));
 OR2_X1 _26238_ (.A1(_02924_),
    .A2(_02960_),
    .ZN(_02970_));
 AOI21_X1 _26239_ (.A(_02747_),
    .B1(_02907_),
    .B2(_02866_),
    .ZN(_02971_));
 AOI21_X1 _26240_ (.A(_02971_),
    .B1(_02937_),
    .B2(_02907_),
    .ZN(_02972_));
 INV_X1 _26241_ (.A(_02972_),
    .ZN(_02973_));
 AOI21_X1 _26242_ (.A(_02903_),
    .B1(_21840_),
    .B2(_02973_),
    .ZN(_02974_));
 AOI21_X1 _26243_ (.A(_02868_),
    .B1(_02835_),
    .B2(_02876_),
    .ZN(_02975_));
 NOR3_X1 _26244_ (.A1(_02908_),
    .A2(_02783_),
    .A3(_02911_),
    .ZN(_02976_));
 OR4_X1 _26245_ (.A1(_02899_),
    .A2(_21840_),
    .A3(_02975_),
    .A4(_02976_),
    .ZN(_02977_));
 AOI221_X2 _26246_ (.A(_02968_),
    .B1(_02969_),
    .B2(_02970_),
    .C1(_02974_),
    .C2(_02977_),
    .ZN(_02978_));
 INV_X2 _26247_ (.A(_02856_),
    .ZN(_02979_));
 MUX2_X1 _26248_ (.A(_02899_),
    .B(_02896_),
    .S(_02979_),
    .Z(_02980_));
 NOR3_X4 _26249_ (.A1(_02961_),
    .A2(_02978_),
    .A3(_02980_),
    .ZN(_02981_));
 XNOR2_X2 _26250_ (.A(_21819_),
    .B(_02840_),
    .ZN(_02982_));
 OAI21_X1 _26251_ (.A(_02922_),
    .B1(_02923_),
    .B2(_02835_),
    .ZN(_02983_));
 NAND2_X1 _26252_ (.A1(_02882_),
    .A2(_02827_),
    .ZN(_02984_));
 AOI21_X1 _26253_ (.A(_02984_),
    .B1(_02835_),
    .B2(_02876_),
    .ZN(_02985_));
 NOR4_X1 _26254_ (.A1(_02905_),
    .A2(_02908_),
    .A3(_02911_),
    .A4(_02902_),
    .ZN(_02986_));
 AOI21_X1 _26255_ (.A(_02903_),
    .B1(_02892_),
    .B2(_02884_),
    .ZN(_02987_));
 OR3_X1 _26256_ (.A1(_02985_),
    .A2(_02986_),
    .A3(_02987_),
    .ZN(_02988_));
 NAND2_X1 _26257_ (.A1(_02983_),
    .A2(_02988_),
    .ZN(_02989_));
 MUX2_X1 _26258_ (.A(_02933_),
    .B(_02939_),
    .S(_02906_),
    .Z(_02990_));
 NAND3_X2 _26259_ (.A1(_02982_),
    .A2(_02989_),
    .A3(_02990_),
    .ZN(_02991_));
 MUX2_X1 _26260_ (.A(_02775_),
    .B(_02783_),
    .S(_02906_),
    .Z(_02992_));
 NAND2_X1 _26261_ (.A1(_02903_),
    .A2(_02868_),
    .ZN(_02993_));
 OAI21_X1 _26262_ (.A(_02993_),
    .B1(_02804_),
    .B2(_02903_),
    .ZN(_02994_));
 MUX2_X1 _26263_ (.A(_02992_),
    .B(_02994_),
    .S(_02940_),
    .Z(_02995_));
 NOR2_X1 _26264_ (.A1(_02995_),
    .A2(_02982_),
    .ZN(_02996_));
 NOR2_X2 _26265_ (.A1(_02855_),
    .A2(_02996_),
    .ZN(_02997_));
 MUX2_X1 _26266_ (.A(_02866_),
    .B(_02896_),
    .S(_02920_),
    .Z(_02998_));
 AOI22_X4 _26267_ (.A1(_02991_),
    .A2(_02997_),
    .B1(_02998_),
    .B2(_02855_),
    .ZN(_02999_));
 AOI21_X1 _26268_ (.A(_02921_),
    .B1(_02869_),
    .B2(_02979_),
    .ZN(_03000_));
 NOR3_X2 _26269_ (.A1(_02855_),
    .A2(_02873_),
    .A3(_02874_),
    .ZN(_03001_));
 AND3_X1 _26270_ (.A1(_02876_),
    .A2(_02800_),
    .A3(_02879_),
    .ZN(_03002_));
 NOR2_X2 _26271_ (.A1(_03001_),
    .A2(_03002_),
    .ZN(_03003_));
 NOR2_X1 _26272_ (.A1(_02852_),
    .A2(_03003_),
    .ZN(_03004_));
 AOI221_X2 _26273_ (.A(_03000_),
    .B1(_03004_),
    .B2(_02988_),
    .C1(_02995_),
    .C2(_02881_),
    .ZN(_03005_));
 NOR2_X2 _26274_ (.A1(_02979_),
    .A2(_02921_),
    .ZN(_03006_));
 AOI21_X4 _26275_ (.A(_03005_),
    .B1(_03006_),
    .B2(_02838_),
    .ZN(_03007_));
 OR2_X1 _26276_ (.A1(_02770_),
    .A2(_02771_),
    .ZN(_03008_));
 NAND2_X1 _26277_ (.A1(_02920_),
    .A2(_03008_),
    .ZN(_03009_));
 OAI221_X2 _26278_ (.A(_03009_),
    .B1(_02896_),
    .B2(_02899_),
    .C1(_02920_),
    .C2(_02798_),
    .ZN(_03010_));
 BUF_X4 _26279_ (.A(_02921_),
    .Z(_03011_));
 NAND4_X2 _26280_ (.A1(_21817_),
    .A2(_03011_),
    .A3(_02924_),
    .A4(_02982_),
    .ZN(_03012_));
 INV_X2 _26281_ (.A(_21819_),
    .ZN(_03013_));
 NOR3_X1 _26282_ (.A1(_02763_),
    .A2(_02764_),
    .A3(_02839_),
    .ZN(_03014_));
 NOR2_X1 _26283_ (.A1(_03013_),
    .A2(_03014_),
    .ZN(_03015_));
 AOI21_X1 _26284_ (.A(_03015_),
    .B1(_02840_),
    .B2(_03013_),
    .ZN(_03016_));
 NOR2_X1 _26285_ (.A1(_02855_),
    .A2(_03016_),
    .ZN(_03017_));
 INV_X1 _26286_ (.A(_02872_),
    .ZN(_03018_));
 NAND2_X1 _26287_ (.A1(_03014_),
    .A2(_03018_),
    .ZN(_03019_));
 OAI21_X2 _26288_ (.A(_03017_),
    .B1(_03019_),
    .B2(_02953_),
    .ZN(_03020_));
 NOR2_X2 _26289_ (.A1(_02903_),
    .A2(_03020_),
    .ZN(_03021_));
 NOR2_X1 _26290_ (.A1(_02906_),
    .A2(_03020_),
    .ZN(_03022_));
 AOI22_X4 _26291_ (.A1(_02950_),
    .A2(_03021_),
    .B1(_03022_),
    .B2(_02955_),
    .ZN(_03023_));
 OAI21_X1 _26292_ (.A(_21840_),
    .B1(_03001_),
    .B2(_03002_),
    .ZN(_03024_));
 NOR4_X1 _26293_ (.A1(_02903_),
    .A2(_03024_),
    .A3(_02975_),
    .A4(_02976_),
    .ZN(_03025_));
 NOR3_X1 _26294_ (.A1(_02906_),
    .A2(_03024_),
    .A3(_02966_),
    .ZN(_03026_));
 NOR2_X1 _26295_ (.A1(_03025_),
    .A2(_03026_),
    .ZN(_03027_));
 NAND4_X4 _26296_ (.A1(_03010_),
    .A2(_03012_),
    .A3(_03023_),
    .A4(_03027_),
    .ZN(_03028_));
 XNOR2_X2 _26297_ (.A(_03013_),
    .B(_02840_),
    .ZN(_03029_));
 NOR4_X2 _26298_ (.A1(_02855_),
    .A2(_02942_),
    .A3(_02943_),
    .A4(_03029_),
    .ZN(_03030_));
 NAND2_X1 _26299_ (.A1(_02921_),
    .A2(_03029_),
    .ZN(_03031_));
 AND2_X1 _26300_ (.A1(_02921_),
    .A2(_02874_),
    .ZN(_03032_));
 OAI221_X1 _26301_ (.A(_02927_),
    .B1(_03019_),
    .B2(_02855_),
    .C1(_02908_),
    .C2(_02911_),
    .ZN(_03033_));
 AOI21_X1 _26302_ (.A(_03032_),
    .B1(_02931_),
    .B2(_03033_),
    .ZN(_03034_));
 MUX2_X1 _26303_ (.A(_02748_),
    .B(_02937_),
    .S(_02979_),
    .Z(_03035_));
 OAI22_X2 _26304_ (.A1(_03031_),
    .A2(_03034_),
    .B1(_03035_),
    .B2(_03011_),
    .ZN(_03036_));
 NOR2_X2 _26305_ (.A1(_03030_),
    .A2(_03036_),
    .ZN(_03037_));
 NAND2_X1 _26306_ (.A1(_02979_),
    .A2(_02747_),
    .ZN(_03038_));
 OAI221_X2 _26307_ (.A(_03038_),
    .B1(_02896_),
    .B2(_02899_),
    .C1(_02979_),
    .C2(_02866_),
    .ZN(_03039_));
 INV_X1 _26308_ (.A(_02783_),
    .ZN(_03040_));
 NOR3_X1 _26309_ (.A1(_03040_),
    .A2(_02951_),
    .A3(_02883_),
    .ZN(_03041_));
 AOI21_X1 _26310_ (.A(_02947_),
    .B1(_02951_),
    .B2(_02804_),
    .ZN(_03042_));
 OAI21_X1 _26311_ (.A(_02886_),
    .B1(_02953_),
    .B2(_02804_),
    .ZN(_03043_));
 NOR2_X1 _26312_ (.A1(_02792_),
    .A2(_02883_),
    .ZN(_03044_));
 AOI221_X2 _26313_ (.A(_03041_),
    .B1(_03042_),
    .B2(_03043_),
    .C1(_03044_),
    .C2(_02836_),
    .ZN(_03045_));
 AND2_X1 _26314_ (.A1(_02851_),
    .A2(_03045_),
    .ZN(_03046_));
 NAND2_X1 _26315_ (.A1(_02875_),
    .A2(_02880_),
    .ZN(_03047_));
 OAI221_X1 _26316_ (.A(_21840_),
    .B1(_02947_),
    .B2(_02966_),
    .C1(_02972_),
    .C2(_02883_),
    .ZN(_03048_));
 NAND2_X1 _26317_ (.A1(_03047_),
    .A2(_03048_),
    .ZN(_03049_));
 NOR4_X2 _26318_ (.A1(_03013_),
    .A2(_02837_),
    .A3(_02867_),
    .A4(_02923_),
    .ZN(_03050_));
 AOI22_X2 _26319_ (.A1(_03013_),
    .A2(_03032_),
    .B1(_03050_),
    .B2(_21816_),
    .ZN(_03051_));
 NOR2_X1 _26320_ (.A1(_02904_),
    .A2(_02912_),
    .ZN(_03052_));
 OAI221_X2 _26321_ (.A(_03039_),
    .B1(_03046_),
    .B2(_03049_),
    .C1(_03051_),
    .C2(_03052_),
    .ZN(_03053_));
 NAND4_X4 _26322_ (.A1(_03007_),
    .A2(_03028_),
    .A3(_03037_),
    .A4(_03053_),
    .ZN(_03054_));
 AOI21_X1 _26323_ (.A(_02921_),
    .B1(_02886_),
    .B2(_02979_),
    .ZN(_03055_));
 NOR4_X1 _26324_ (.A1(_02985_),
    .A2(_02986_),
    .A3(_02987_),
    .A4(_03055_),
    .ZN(_03056_));
 NAND2_X1 _26325_ (.A1(_02804_),
    .A2(_03006_),
    .ZN(_03057_));
 OAI21_X1 _26326_ (.A(_03057_),
    .B1(_03055_),
    .B2(_02881_),
    .ZN(_03058_));
 NOR2_X1 _26327_ (.A1(_03056_),
    .A2(_03058_),
    .ZN(_21822_));
 AND2_X1 _26328_ (.A1(_21821_),
    .A2(_21822_),
    .ZN(_03059_));
 NOR2_X1 _26329_ (.A1(_02979_),
    .A2(_02868_),
    .ZN(_03060_));
 NOR2_X1 _26330_ (.A1(_02920_),
    .A2(_02783_),
    .ZN(_03061_));
 NOR2_X1 _26331_ (.A1(_21840_),
    .A2(_02893_),
    .ZN(_03062_));
 AND3_X1 _26332_ (.A1(_21840_),
    .A2(_02928_),
    .A3(_02931_),
    .ZN(_03063_));
 OAI33_X1 _26333_ (.A1(_02921_),
    .A2(_03060_),
    .A3(_03061_),
    .B1(_03062_),
    .B2(_03063_),
    .B3(_03003_),
    .ZN(_03064_));
 NOR2_X1 _26334_ (.A1(_02856_),
    .A2(_02804_),
    .ZN(_03065_));
 AOI21_X2 _26335_ (.A(_03065_),
    .B1(_02783_),
    .B2(_02920_),
    .ZN(_03066_));
 OAI22_X4 _26336_ (.A1(_03003_),
    .A2(_02957_),
    .B1(_03066_),
    .B2(_02921_),
    .ZN(_03067_));
 OAI21_X1 _26337_ (.A(_02855_),
    .B1(_02868_),
    .B2(_02856_),
    .ZN(_03068_));
 OAI21_X1 _26338_ (.A(_02711_),
    .B1(_02904_),
    .B2(_02912_),
    .ZN(_03069_));
 OAI221_X1 _26339_ (.A(_03068_),
    .B1(_03020_),
    .B2(_03069_),
    .C1(_03024_),
    .C2(_03045_),
    .ZN(_03070_));
 NAND2_X1 _26340_ (.A1(_02869_),
    .A2(_03006_),
    .ZN(_03071_));
 AND2_X2 _26341_ (.A1(_03070_),
    .A2(_03071_),
    .ZN(_03072_));
 NAND4_X4 _26342_ (.A1(_03059_),
    .A2(_03064_),
    .A3(_03067_),
    .A4(_03072_),
    .ZN(_03073_));
 NOR4_X4 _26343_ (.A1(_02981_),
    .A2(_02999_),
    .A3(_03054_),
    .A4(_03073_),
    .ZN(_03074_));
 XOR2_X1 _26344_ (.A(_02946_),
    .B(_03074_),
    .Z(_03075_));
 AND2_X1 _26345_ (.A1(_21824_),
    .A2(_03075_),
    .ZN(_03076_));
 BUF_X4 _26346_ (.A(_03075_),
    .Z(_21827_));
 NAND2_X1 _26347_ (.A1(_02893_),
    .A2(_03069_),
    .ZN(_03077_));
 NAND3_X1 _26348_ (.A1(_21817_),
    .A2(_21840_),
    .A3(_21844_),
    .ZN(_03078_));
 AOI21_X1 _26349_ (.A(_03077_),
    .B1(_03078_),
    .B2(_03011_),
    .ZN(_03079_));
 NOR2_X1 _26350_ (.A1(_02893_),
    .A2(_03069_),
    .ZN(_03080_));
 OAI21_X1 _26351_ (.A(_02881_),
    .B1(_03079_),
    .B2(_03080_),
    .ZN(_03081_));
 XNOR2_X1 _26352_ (.A(_02865_),
    .B(_02900_),
    .ZN(_03082_));
 AOI21_X1 _26353_ (.A(_21827_),
    .B1(_03081_),
    .B2(_03082_),
    .ZN(_03083_));
 NOR3_X1 _26354_ (.A1(_02491_),
    .A2(_03076_),
    .A3(_03083_),
    .ZN(_03084_));
 OAI21_X1 _26355_ (.A(_02915_),
    .B1(_02919_),
    .B2(_03084_),
    .ZN(_00096_));
 NAND2_X1 _26356_ (.A1(\g_reduce0[6].adder.b[1] ),
    .A2(_02914_),
    .ZN(_03085_));
 XOR2_X2 _26357_ (.A(_21823_),
    .B(_03067_),
    .Z(_03086_));
 NOR2_X1 _26358_ (.A1(_02491_),
    .A2(_03086_),
    .ZN(_03087_));
 NAND2_X1 _26359_ (.A1(_21827_),
    .A2(_03087_),
    .ZN(_03088_));
 OR2_X1 _26360_ (.A1(_21824_),
    .A2(_02491_),
    .ZN(_03089_));
 OAI221_X2 _26361_ (.A(_03088_),
    .B1(_03089_),
    .B2(_21827_),
    .C1(\g_reduce0[6].adder.a[1] ),
    .C2(_02918_),
    .ZN(_03090_));
 OAI21_X1 _26362_ (.A(_03085_),
    .B1(_03090_),
    .B2(_02914_),
    .ZN(_00103_));
 NOR2_X1 _26363_ (.A1(\g_reduce0[6].adder.a[2] ),
    .A2(_02918_),
    .ZN(_03091_));
 NOR3_X1 _26364_ (.A1(_02491_),
    .A2(_03075_),
    .A3(_03086_),
    .ZN(_03092_));
 NAND2_X1 _26365_ (.A1(_03059_),
    .A2(_03067_),
    .ZN(_03093_));
 XOR2_X2 _26366_ (.A(net341),
    .B(_03093_),
    .Z(_03094_));
 AND3_X1 _26367_ (.A1(_02918_),
    .A2(_03075_),
    .A3(_03094_),
    .ZN(_03095_));
 NOR3_X1 _26368_ (.A1(_03091_),
    .A2(_03092_),
    .A3(_03095_),
    .ZN(_03096_));
 MUX2_X1 _26369_ (.A(\g_reduce0[6].adder.b[2] ),
    .B(_03096_),
    .S(_02916_),
    .Z(_00104_));
 NOR2_X1 _26370_ (.A1(\g_reduce0[6].adder.b[3] ),
    .A2(_02916_),
    .ZN(_03097_));
 AOI21_X1 _26371_ (.A(_02914_),
    .B1(_02491_),
    .B2(\g_reduce0[6].adder.a[3] ),
    .ZN(_03098_));
 NAND3_X1 _26372_ (.A1(_21823_),
    .A2(net341),
    .A3(_03067_),
    .ZN(_03099_));
 XOR2_X2 _26373_ (.A(_03072_),
    .B(_03099_),
    .Z(_03100_));
 MUX2_X1 _26374_ (.A(_03094_),
    .B(_03100_),
    .S(_03075_),
    .Z(_03101_));
 OR2_X1 _26375_ (.A1(_02491_),
    .A2(_03101_),
    .ZN(_03102_));
 AOI21_X1 _26376_ (.A(_03097_),
    .B1(_03098_),
    .B2(_03102_),
    .ZN(_00105_));
 NOR2_X1 _26377_ (.A1(_02914_),
    .A2(_02918_),
    .ZN(_03103_));
 AOI22_X1 _26378_ (.A1(\g_reduce0[6].adder.b[4] ),
    .A2(_02914_),
    .B1(_03103_),
    .B2(\g_reduce0[6].adder.a[4] ),
    .ZN(_03104_));
 XOR2_X2 _26379_ (.A(_03007_),
    .B(_03073_),
    .Z(_03105_));
 MUX2_X1 _26380_ (.A(_03100_),
    .B(_03105_),
    .S(_21827_),
    .Z(_03106_));
 NAND2_X1 _26381_ (.A1(_02486_),
    .A2(_02917_),
    .ZN(_03107_));
 OAI21_X1 _26382_ (.A(_03104_),
    .B1(_03106_),
    .B2(_03107_),
    .ZN(_00106_));
 NOR2_X2 _26383_ (.A1(_02914_),
    .A2(_02491_),
    .ZN(_03108_));
 AND4_X1 _26384_ (.A1(_21823_),
    .A2(net341),
    .A3(_03067_),
    .A4(_03072_),
    .ZN(_03109_));
 NAND2_X1 _26385_ (.A1(_03007_),
    .A2(_03109_),
    .ZN(_03110_));
 XOR2_X2 _26386_ (.A(_03028_),
    .B(_03110_),
    .Z(_03111_));
 AND3_X1 _26387_ (.A1(_21827_),
    .A2(_03108_),
    .A3(_03111_),
    .ZN(_03112_));
 NAND2_X1 _26388_ (.A1(_03108_),
    .A2(_03105_),
    .ZN(_03113_));
 NOR2_X1 _26389_ (.A1(_21827_),
    .A2(_03113_),
    .ZN(_03114_));
 NAND2_X1 _26390_ (.A1(_02486_),
    .A2(_02491_),
    .ZN(_03115_));
 OAI22_X1 _26391_ (.A1(\g_reduce0[6].adder.b[5] ),
    .A2(_02916_),
    .B1(_03115_),
    .B2(\g_reduce0[6].adder.a[5] ),
    .ZN(_03116_));
 NOR3_X1 _26392_ (.A1(_03112_),
    .A2(_03114_),
    .A3(_03116_),
    .ZN(_00107_));
 NAND2_X1 _26393_ (.A1(_03108_),
    .A2(_03111_),
    .ZN(_03117_));
 NOR2_X1 _26394_ (.A1(_21827_),
    .A2(_03117_),
    .ZN(_03118_));
 INV_X1 _26395_ (.A(_03073_),
    .ZN(_03119_));
 AND3_X1 _26396_ (.A1(_03007_),
    .A2(_03028_),
    .A3(_03119_),
    .ZN(_03120_));
 XNOR2_X1 _26397_ (.A(_03037_),
    .B(_03120_),
    .ZN(_03121_));
 AND3_X1 _26398_ (.A1(_21827_),
    .A2(_03108_),
    .A3(_03121_),
    .ZN(_03122_));
 OAI22_X1 _26399_ (.A1(\g_reduce0[6].adder.b[6] ),
    .A2(_02916_),
    .B1(_03115_),
    .B2(\g_reduce0[6].adder.a[6] ),
    .ZN(_03123_));
 NOR3_X1 _26400_ (.A1(_03118_),
    .A2(_03122_),
    .A3(_03123_),
    .ZN(_00108_));
 OAI22_X1 _26401_ (.A1(\g_reduce0[6].adder.b[7] ),
    .A2(_02916_),
    .B1(_03115_),
    .B2(\g_reduce0[6].adder.a[7] ),
    .ZN(_03124_));
 NAND4_X1 _26402_ (.A1(_03007_),
    .A2(_03028_),
    .A3(_03037_),
    .A4(_03109_),
    .ZN(_03125_));
 XOR2_X2 _26403_ (.A(_03053_),
    .B(_03125_),
    .Z(_03126_));
 MUX2_X1 _26404_ (.A(_03121_),
    .B(_03126_),
    .S(_21827_),
    .Z(_03127_));
 AOI21_X1 _26405_ (.A(_03124_),
    .B1(_03127_),
    .B2(_03108_),
    .ZN(_00109_));
 OAI21_X1 _26406_ (.A(_02999_),
    .B1(_03054_),
    .B2(_03073_),
    .ZN(_03128_));
 NOR2_X1 _26407_ (.A1(_02981_),
    .A2(_03109_),
    .ZN(_03129_));
 OR3_X1 _26408_ (.A1(_02999_),
    .A2(_03054_),
    .A3(_03073_),
    .ZN(_03130_));
 OAI21_X1 _26409_ (.A(_03128_),
    .B1(_03129_),
    .B2(_03130_),
    .ZN(_03131_));
 NAND2_X1 _26410_ (.A1(_02946_),
    .A2(_03108_),
    .ZN(_03132_));
 NOR2_X1 _26411_ (.A1(_03131_),
    .A2(_03132_),
    .ZN(_03133_));
 NOR2_X1 _26412_ (.A1(_02946_),
    .A2(_03107_),
    .ZN(_03134_));
 NOR2_X1 _26413_ (.A1(_03074_),
    .A2(_03126_),
    .ZN(_03135_));
 AOI21_X1 _26414_ (.A(_03133_),
    .B1(_03134_),
    .B2(_03135_),
    .ZN(_03136_));
 AOI22_X1 _26415_ (.A1(\g_reduce0[6].adder.b[8] ),
    .A2(_02914_),
    .B1(_03103_),
    .B2(\g_reduce0[6].adder.a[8] ),
    .ZN(_03137_));
 NAND2_X1 _26416_ (.A1(_03136_),
    .A2(_03137_),
    .ZN(_00110_));
 NAND2_X1 _26417_ (.A1(_03131_),
    .A2(_03134_),
    .ZN(_03138_));
 NOR2_X1 _26418_ (.A1(_02999_),
    .A2(_03054_),
    .ZN(_03139_));
 OAI21_X1 _26419_ (.A(_03139_),
    .B1(_03119_),
    .B2(_03109_),
    .ZN(_03140_));
 AND2_X1 _26420_ (.A1(_03139_),
    .A2(_03109_),
    .ZN(_03141_));
 MUX2_X1 _26421_ (.A(_03140_),
    .B(_03141_),
    .S(_02981_),
    .Z(_03142_));
 OAI221_X1 _26422_ (.A(_03138_),
    .B1(_03142_),
    .B2(_03132_),
    .C1(_03115_),
    .C2(\g_reduce0[6].adder.a[9] ),
    .ZN(_03143_));
 INV_X1 _26423_ (.A(\g_reduce0[6].adder.b[9] ),
    .ZN(_03144_));
 AOI21_X1 _26424_ (.A(_03143_),
    .B1(_02914_),
    .B2(_03144_),
    .ZN(_00111_));
 INV_X1 _26425_ (.A(_21825_),
    .ZN(_21831_));
 MUX2_X1 _26426_ (.A(\g_reduce0[6].adder.a[10] ),
    .B(_21830_),
    .S(_02918_),
    .Z(_03145_));
 MUX2_X1 _26427_ (.A(\g_reduce0[6].adder.b[10] ),
    .B(_03145_),
    .S(_02916_),
    .Z(_00097_));
 MUX2_X1 _26428_ (.A(_02482_),
    .B(_21838_),
    .S(_02918_),
    .Z(_03146_));
 MUX2_X1 _26429_ (.A(_02487_),
    .B(_03146_),
    .S(_02916_),
    .Z(_00098_));
 MUX2_X2 _26430_ (.A(_21703_),
    .B(_00542_),
    .S(_02532_),
    .Z(_03147_));
 NAND2_X1 _26431_ (.A1(_02920_),
    .A2(_21832_),
    .ZN(_03148_));
 XOR2_X1 _26432_ (.A(_03147_),
    .B(_03148_),
    .Z(_03149_));
 XOR2_X1 _26433_ (.A(_14130_),
    .B(_21842_),
    .Z(_03150_));
 MUX2_X1 _26434_ (.A(_03149_),
    .B(_03150_),
    .S(_03011_),
    .Z(_03151_));
 XOR2_X1 _26435_ (.A(_21837_),
    .B(_03151_),
    .Z(_03152_));
 MUX2_X1 _26436_ (.A(_02483_),
    .B(_03152_),
    .S(_02918_),
    .Z(_03153_));
 MUX2_X1 _26437_ (.A(_02488_),
    .B(_03153_),
    .S(_02916_),
    .Z(_00099_));
 INV_X1 _26438_ (.A(_14132_),
    .ZN(_14129_));
 MUX2_X1 _26439_ (.A(_21700_),
    .B(_00545_),
    .S(_02533_),
    .Z(_03154_));
 MUX2_X1 _26440_ (.A(_21706_),
    .B(_00537_),
    .S(_02533_),
    .Z(_03155_));
 NOR4_X1 _26441_ (.A1(_02979_),
    .A2(_21825_),
    .A3(_03147_),
    .A4(_03155_),
    .ZN(_03156_));
 XNOR2_X1 _26442_ (.A(_03154_),
    .B(_03156_),
    .ZN(_03157_));
 INV_X1 _26443_ (.A(_21834_),
    .ZN(_03158_));
 INV_X1 _26444_ (.A(_21835_),
    .ZN(_03159_));
 OAI21_X1 _26445_ (.A(_03158_),
    .B1(_03159_),
    .B2(_14132_),
    .ZN(_03160_));
 AOI21_X1 _26446_ (.A(_21841_),
    .B1(_03160_),
    .B2(_21842_),
    .ZN(_03161_));
 XNOR2_X1 _26447_ (.A(_21846_),
    .B(_03161_),
    .ZN(_03162_));
 MUX2_X1 _26448_ (.A(_03157_),
    .B(_03162_),
    .S(_03011_),
    .Z(_03163_));
 NAND2_X1 _26449_ (.A1(_02920_),
    .A2(_21833_),
    .ZN(_03164_));
 OAI21_X1 _26450_ (.A(_03164_),
    .B1(_03155_),
    .B2(_02920_),
    .ZN(_03165_));
 MUX2_X1 _26451_ (.A(_14131_),
    .B(_03165_),
    .S(_02855_),
    .Z(_21836_));
 NAND3_X1 _26452_ (.A1(_21829_),
    .A2(_03151_),
    .A3(_21836_),
    .ZN(_03166_));
 XNOR2_X1 _26453_ (.A(_03163_),
    .B(_03166_),
    .ZN(_03167_));
 MUX2_X1 _26454_ (.A(\g_reduce0[6].adder.a[13] ),
    .B(_03167_),
    .S(_02918_),
    .Z(_03168_));
 MUX2_X1 _26455_ (.A(\g_reduce0[6].adder.b[13] ),
    .B(_03168_),
    .S(_02916_),
    .Z(_00100_));
 INV_X1 _26456_ (.A(_02489_),
    .ZN(_03169_));
 NOR2_X1 _26457_ (.A1(_03169_),
    .A2(_02545_),
    .ZN(_03170_));
 NOR2_X1 _26458_ (.A1(_02489_),
    .A2(_02486_),
    .ZN(_03171_));
 NOR3_X1 _26459_ (.A1(_02484_),
    .A2(_03170_),
    .A3(_03171_),
    .ZN(_03172_));
 NOR4_X1 _26460_ (.A1(_03011_),
    .A2(_03147_),
    .A3(_03148_),
    .A4(_03154_),
    .ZN(_03173_));
 AOI21_X1 _26461_ (.A(_21841_),
    .B1(_21842_),
    .B2(_14130_),
    .ZN(_03174_));
 INV_X1 _26462_ (.A(_03174_),
    .ZN(_03175_));
 AOI21_X1 _26463_ (.A(_21845_),
    .B1(_03175_),
    .B2(_21846_),
    .ZN(_03176_));
 AOI21_X1 _26464_ (.A(_03173_),
    .B1(_03176_),
    .B2(_03011_),
    .ZN(_03177_));
 NAND3_X1 _26465_ (.A1(_21837_),
    .A2(_03151_),
    .A3(_03163_),
    .ZN(_03178_));
 XNOR2_X2 _26466_ (.A(_03177_),
    .B(_03178_),
    .ZN(_03179_));
 MUX2_X1 _26467_ (.A(_03172_),
    .B(_03170_),
    .S(_03179_),
    .Z(_03180_));
 AOI21_X1 _26468_ (.A(_02491_),
    .B1(_02545_),
    .B2(_03179_),
    .ZN(_03181_));
 NAND2_X1 _26469_ (.A1(_03169_),
    .A2(_02505_),
    .ZN(_03182_));
 OAI21_X1 _26470_ (.A(_03181_),
    .B1(_03182_),
    .B2(_03179_),
    .ZN(_03183_));
 AOI222_X2 _26471_ (.A1(_02489_),
    .A2(_02914_),
    .B1(_02918_),
    .B2(_03180_),
    .C1(_03183_),
    .C2(_02484_),
    .ZN(_03184_));
 INV_X1 _26472_ (.A(_03184_),
    .ZN(_00101_));
 BUF_X2 _26473_ (.A(\g_reduce0[8].adder.a[11] ),
    .Z(_03185_));
 CLKBUF_X2 _26474_ (.A(\g_reduce0[8].adder.a[10] ),
    .Z(_03186_));
 OR2_X1 _26475_ (.A1(_03186_),
    .A2(\g_reduce0[8].adder.a[13] ),
    .ZN(_03187_));
 OR4_X1 _26476_ (.A1(_03185_),
    .A2(\g_reduce0[8].adder.a[12] ),
    .A3(\g_reduce0[8].adder.a[14] ),
    .A4(_03187_),
    .ZN(_03188_));
 CLKBUF_X3 _26477_ (.A(_03188_),
    .Z(_03189_));
 BUF_X2 _26478_ (.A(\g_reduce0[8].adder.b[14] ),
    .Z(_03190_));
 OR2_X1 _26479_ (.A1(\g_reduce0[8].adder.b[10] ),
    .A2(\g_reduce0[8].adder.b[13] ),
    .ZN(_03191_));
 NOR4_X4 _26480_ (.A1(\g_reduce0[8].adder.b[11] ),
    .A2(\g_reduce0[8].adder.b[12] ),
    .A3(_03190_),
    .A4(_03191_),
    .ZN(_03192_));
 INV_X1 _26481_ (.A(_21890_),
    .ZN(_03193_));
 INV_X1 _26482_ (.A(_21851_),
    .ZN(_03194_));
 INV_X1 _26483_ (.A(_21857_),
    .ZN(_03195_));
 AOI21_X1 _26484_ (.A(_21854_),
    .B1(_03195_),
    .B2(_21855_),
    .ZN(_03196_));
 BUF_X1 _26485_ (.A(_21852_),
    .Z(_03197_));
 INV_X2 _26486_ (.A(_03197_),
    .ZN(_03198_));
 OAI21_X1 _26487_ (.A(_03194_),
    .B1(_03196_),
    .B2(_03198_),
    .ZN(_03199_));
 BUF_X2 _26488_ (.A(_21849_),
    .Z(_03200_));
 AOI21_X2 _26489_ (.A(_21848_),
    .B1(_03199_),
    .B2(_03200_),
    .ZN(_03201_));
 CLKBUF_X3 _26490_ (.A(_21891_),
    .Z(_03202_));
 INV_X4 _26491_ (.A(_03202_),
    .ZN(_03203_));
 OAI21_X4 _26492_ (.A(_03193_),
    .B1(_03201_),
    .B2(_03203_),
    .ZN(_03204_));
 AND4_X1 _26493_ (.A1(_21861_),
    .A2(_21864_),
    .A3(_21867_),
    .A4(_21870_),
    .ZN(_03205_));
 NOR2_X1 _26494_ (.A1(_21881_),
    .A2(_21872_),
    .ZN(_03206_));
 AOI21_X1 _26495_ (.A(_21875_),
    .B1(_21878_),
    .B2(_21876_),
    .ZN(_03207_));
 INV_X1 _26496_ (.A(_21873_),
    .ZN(_03208_));
 OAI21_X1 _26497_ (.A(_03206_),
    .B1(_03207_),
    .B2(_03208_),
    .ZN(_03209_));
 INV_X1 _26498_ (.A(_21882_),
    .ZN(_03210_));
 INV_X1 _26499_ (.A(_21884_),
    .ZN(_03211_));
 INV_X1 _26500_ (.A(\g_reduce0[8].adder.a[0] ),
    .ZN(_03212_));
 OAI21_X1 _26501_ (.A(_21885_),
    .B1(\g_reduce0[8].adder.b[0] ),
    .B2(_03212_),
    .ZN(_03213_));
 AOI21_X1 _26502_ (.A(_03210_),
    .B1(_03211_),
    .B2(_03213_),
    .ZN(_03214_));
 INV_X1 _26503_ (.A(_21875_),
    .ZN(_03215_));
 OAI21_X1 _26504_ (.A(_21876_),
    .B1(_21879_),
    .B2(_21878_),
    .ZN(_03216_));
 AOI21_X1 _26505_ (.A(_03208_),
    .B1(_03215_),
    .B2(_03216_),
    .ZN(_03217_));
 OAI221_X2 _26506_ (.A(_03205_),
    .B1(_03209_),
    .B2(_03214_),
    .C1(_03217_),
    .C2(_21872_),
    .ZN(_03218_));
 INV_X1 _26507_ (.A(_21863_),
    .ZN(_03219_));
 AOI21_X1 _26508_ (.A(_21866_),
    .B1(_21867_),
    .B2(_21869_),
    .ZN(_03220_));
 INV_X1 _26509_ (.A(_21864_),
    .ZN(_03221_));
 OAI21_X1 _26510_ (.A(_03219_),
    .B1(_03220_),
    .B2(_03221_),
    .ZN(_03222_));
 AND2_X1 _26511_ (.A1(_21861_),
    .A2(_03222_),
    .ZN(_03223_));
 CLKBUF_X3 _26512_ (.A(_21858_),
    .Z(_03224_));
 NAND4_X2 _26513_ (.A1(_03224_),
    .A2(_03200_),
    .A3(_03197_),
    .A4(_21855_),
    .ZN(_03225_));
 NOR4_X4 _26514_ (.A1(_03203_),
    .A2(_21860_),
    .A3(_03223_),
    .A4(_03225_),
    .ZN(_03226_));
 NAND2_X4 _26515_ (.A1(_03218_),
    .A2(_03226_),
    .ZN(_03227_));
 NAND2_X4 _26516_ (.A1(_03204_),
    .A2(_03227_),
    .ZN(_03228_));
 OAI21_X1 _26517_ (.A(_03189_),
    .B1(_03192_),
    .B2(_03228_),
    .ZN(_03229_));
 MUX2_X1 _26518_ (.A(\g_reduce0[8].adder.a[15] ),
    .B(\g_reduce0[8].adder.b[15] ),
    .S(_03229_),
    .Z(_00118_));
 INV_X1 _26519_ (.A(_21848_),
    .ZN(_03230_));
 INV_X1 _26520_ (.A(_21854_),
    .ZN(_03231_));
 INV_X1 _26521_ (.A(_21855_),
    .ZN(_03232_));
 OAI21_X1 _26522_ (.A(_03231_),
    .B1(_21857_),
    .B2(_03232_),
    .ZN(_03233_));
 AOI21_X1 _26523_ (.A(_21851_),
    .B1(_03233_),
    .B2(_03197_),
    .ZN(_03234_));
 INV_X1 _26524_ (.A(_03200_),
    .ZN(_03235_));
 OAI21_X2 _26525_ (.A(_03230_),
    .B1(_03234_),
    .B2(_03235_),
    .ZN(_03236_));
 AOI21_X4 _26526_ (.A(_21890_),
    .B1(_03236_),
    .B2(_03202_),
    .ZN(_03237_));
 AND2_X1 _26527_ (.A1(_03218_),
    .A2(_03226_),
    .ZN(_03238_));
 BUF_X4 _26528_ (.A(_03238_),
    .Z(_03239_));
 NOR2_X4 _26529_ (.A1(_03237_),
    .A2(_03239_),
    .ZN(_03240_));
 MUX2_X1 _26530_ (.A(_03186_),
    .B(\g_reduce0[8].adder.b[10] ),
    .S(_03240_),
    .Z(_21975_));
 OR4_X1 _26531_ (.A1(\g_reduce0[8].adder.a[13] ),
    .A2(_00559_),
    .A3(_03237_),
    .A4(_03239_),
    .ZN(_03241_));
 NOR2_X1 _26532_ (.A1(\g_reduce0[8].adder.b[13] ),
    .A2(_21847_),
    .ZN(_03242_));
 OAI21_X1 _26533_ (.A(_03242_),
    .B1(_03239_),
    .B2(_03237_),
    .ZN(_03243_));
 NAND2_X2 _26534_ (.A1(_03241_),
    .A2(_03243_),
    .ZN(_03244_));
 NOR2_X2 _26535_ (.A1(\g_reduce0[8].adder.b[11] ),
    .A2(_21853_),
    .ZN(_03245_));
 NOR2_X2 _26536_ (.A1(_21887_),
    .A2(_03245_),
    .ZN(_03246_));
 OAI222_X2 _26537_ (.A1(\g_reduce0[8].adder.b[12] ),
    .A2(_21850_),
    .B1(_03237_),
    .B2(_03239_),
    .C1(_03246_),
    .C2(_03198_),
    .ZN(_03247_));
 OR2_X1 _26538_ (.A1(\g_reduce0[8].adder.a[12] ),
    .A2(_00556_),
    .ZN(_03248_));
 NOR2_X1 _26539_ (.A1(_03185_),
    .A2(_00551_),
    .ZN(_03249_));
 OAI21_X1 _26540_ (.A(_03197_),
    .B1(_03249_),
    .B2(_21887_),
    .ZN(_03250_));
 NAND4_X2 _26541_ (.A1(_03204_),
    .A2(_03227_),
    .A3(_03248_),
    .A4(_03250_),
    .ZN(_03251_));
 AND3_X1 _26542_ (.A1(_03200_),
    .A2(_03247_),
    .A3(_03251_),
    .ZN(_03252_));
 OAI21_X2 _26543_ (.A(_03202_),
    .B1(_03244_),
    .B2(_03252_),
    .ZN(_03253_));
 AND2_X1 _26544_ (.A1(_03241_),
    .A2(_03243_),
    .ZN(_03254_));
 NAND3_X2 _26545_ (.A1(_03200_),
    .A2(_03247_),
    .A3(_03251_),
    .ZN(_03255_));
 NAND3_X2 _26546_ (.A1(_03203_),
    .A2(_03254_),
    .A3(_03255_),
    .ZN(_03256_));
 NAND2_X2 _26547_ (.A1(_03253_),
    .A2(_03256_),
    .ZN(_03257_));
 OR3_X1 _26548_ (.A1(\g_reduce0[8].adder.b[12] ),
    .A2(_21850_),
    .A3(_03240_),
    .ZN(_03258_));
 INV_X1 _26549_ (.A(\g_reduce0[8].adder.b[10] ),
    .ZN(_03259_));
 AND2_X1 _26550_ (.A1(_03186_),
    .A2(_03259_),
    .ZN(_03260_));
 OAI21_X1 _26551_ (.A(_03260_),
    .B1(_00551_),
    .B2(_03185_),
    .ZN(_03261_));
 NOR2_X1 _26552_ (.A1(_03186_),
    .A2(_03245_),
    .ZN(_03262_));
 OAI21_X1 _26553_ (.A(_03262_),
    .B1(_03239_),
    .B2(_03237_),
    .ZN(_03263_));
 OAI221_X2 _26554_ (.A(_03197_),
    .B1(_03228_),
    .B2(_03261_),
    .C1(_03263_),
    .C2(_03259_),
    .ZN(_03264_));
 NAND3_X1 _26555_ (.A1(_03204_),
    .A2(_03227_),
    .A3(_03249_),
    .ZN(_03265_));
 OAI21_X1 _26556_ (.A(_03245_),
    .B1(_03239_),
    .B2(_03237_),
    .ZN(_03266_));
 AND3_X1 _26557_ (.A1(_03232_),
    .A2(_03265_),
    .A3(_03266_),
    .ZN(_03267_));
 OAI221_X2 _26558_ (.A(_03258_),
    .B1(_03264_),
    .B2(_03267_),
    .C1(_03248_),
    .C2(_03228_),
    .ZN(_03268_));
 XNOR2_X2 _26559_ (.A(_03235_),
    .B(_03268_),
    .ZN(_03269_));
 CLKBUF_X3 _26560_ (.A(_03269_),
    .Z(_03270_));
 MUX2_X1 _26561_ (.A(_00554_),
    .B(_21865_),
    .S(_03240_),
    .Z(_03271_));
 CLKBUF_X3 _26562_ (.A(_03240_),
    .Z(_03272_));
 MUX2_X1 _26563_ (.A(_00555_),
    .B(_21868_),
    .S(_03272_),
    .Z(_03273_));
 CLKBUF_X3 _26564_ (.A(_03224_),
    .Z(_03274_));
 MUX2_X1 _26565_ (.A(_03271_),
    .B(_03273_),
    .S(_03274_),
    .Z(_03275_));
 MUX2_X1 _26566_ (.A(_00552_),
    .B(_21871_),
    .S(_03272_),
    .Z(_03276_));
 MUX2_X1 _26567_ (.A(_00553_),
    .B(_21874_),
    .S(_03272_),
    .Z(_03277_));
 MUX2_X1 _26568_ (.A(_03276_),
    .B(_03277_),
    .S(_03274_),
    .Z(_03278_));
 BUF_X4 _26569_ (.A(_21888_),
    .Z(_03279_));
 INV_X2 _26570_ (.A(_03279_),
    .ZN(_03280_));
 MUX2_X1 _26571_ (.A(_03275_),
    .B(_03278_),
    .S(_03280_),
    .Z(_03281_));
 MUX2_X1 _26572_ (.A(_00550_),
    .B(_21880_),
    .S(_03240_),
    .Z(_03282_));
 MUX2_X1 _26573_ (.A(_00549_),
    .B(_21877_),
    .S(_03272_),
    .Z(_03283_));
 INV_X2 _26574_ (.A(_03224_),
    .ZN(_03284_));
 MUX2_X1 _26575_ (.A(_03282_),
    .B(_03283_),
    .S(_03284_),
    .Z(_03285_));
 MUX2_X1 _26576_ (.A(_00546_),
    .B(_21883_),
    .S(_03240_),
    .Z(_03286_));
 MUX2_X1 _26577_ (.A(_00547_),
    .B(_00548_),
    .S(_03272_),
    .Z(_03287_));
 MUX2_X1 _26578_ (.A(_03286_),
    .B(_03287_),
    .S(_03274_),
    .Z(_03288_));
 MUX2_X1 _26579_ (.A(_03285_),
    .B(_03288_),
    .S(_03280_),
    .Z(_03289_));
 OAI21_X2 _26580_ (.A(_03246_),
    .B1(_03239_),
    .B2(_03237_),
    .ZN(_03290_));
 NOR2_X1 _26581_ (.A1(_21887_),
    .A2(_03249_),
    .ZN(_03291_));
 NAND3_X2 _26582_ (.A1(_03204_),
    .A2(_03227_),
    .A3(_03291_),
    .ZN(_03292_));
 NAND3_X1 _26583_ (.A1(_03197_),
    .A2(_03290_),
    .A3(_03292_),
    .ZN(_03293_));
 INV_X1 _26584_ (.A(_03246_),
    .ZN(_03294_));
 AOI21_X2 _26585_ (.A(_03294_),
    .B1(_03227_),
    .B2(_03204_),
    .ZN(_03295_));
 AND3_X1 _26586_ (.A1(_03204_),
    .A2(_03227_),
    .A3(_03291_),
    .ZN(_03296_));
 OAI21_X1 _26587_ (.A(_03198_),
    .B1(_03295_),
    .B2(_03296_),
    .ZN(_03297_));
 NAND2_X2 _26588_ (.A1(_03293_),
    .A2(_03297_),
    .ZN(_03298_));
 CLKBUF_X3 _26589_ (.A(_03298_),
    .Z(_03299_));
 MUX2_X1 _26590_ (.A(_03281_),
    .B(_03289_),
    .S(_03299_),
    .Z(_03300_));
 MUX2_X1 _26591_ (.A(_00558_),
    .B(_21862_),
    .S(_03240_),
    .Z(_03301_));
 MUX2_X1 _26592_ (.A(_00557_),
    .B(_21859_),
    .S(_03272_),
    .Z(_03302_));
 MUX2_X1 _26593_ (.A(_03301_),
    .B(_03302_),
    .S(_03284_),
    .Z(_03303_));
 MUX2_X1 _26594_ (.A(_03284_),
    .B(_03303_),
    .S(_03280_),
    .Z(_03304_));
 NAND2_X1 _26595_ (.A1(_03270_),
    .A2(_03299_),
    .ZN(_03305_));
 OAI22_X1 _26596_ (.A1(_03270_),
    .A2(_03300_),
    .B1(_03304_),
    .B2(_03305_),
    .ZN(_03306_));
 NAND2_X1 _26597_ (.A1(_03257_),
    .A2(_03306_),
    .ZN(_21955_));
 INV_X1 _26598_ (.A(_21955_),
    .ZN(_21952_));
 AOI21_X4 _26599_ (.A(_03203_),
    .B1(_03254_),
    .B2(_03255_),
    .ZN(_03307_));
 NOR3_X4 _26600_ (.A1(_03202_),
    .A2(_03244_),
    .A3(_03252_),
    .ZN(_03308_));
 NOR2_X4 _26601_ (.A1(_03307_),
    .A2(_03308_),
    .ZN(_03309_));
 AND2_X1 _26602_ (.A1(_03224_),
    .A2(_00552_),
    .ZN(_03310_));
 AOI221_X2 _26603_ (.A(_03310_),
    .B1(_03227_),
    .B2(_03204_),
    .C1(_03284_),
    .C2(_00555_),
    .ZN(_03311_));
 MUX2_X1 _26604_ (.A(_21868_),
    .B(_21871_),
    .S(_03224_),
    .Z(_03312_));
 NOR3_X1 _26605_ (.A1(_03237_),
    .A2(_03239_),
    .A3(_03312_),
    .ZN(_03313_));
 NOR2_X1 _26606_ (.A1(_03311_),
    .A2(_03313_),
    .ZN(_03314_));
 MUX2_X1 _26607_ (.A(_03271_),
    .B(_03301_),
    .S(_03284_),
    .Z(_03315_));
 MUX2_X1 _26608_ (.A(_03314_),
    .B(_03315_),
    .S(_03279_),
    .Z(_03316_));
 MUX2_X1 _26609_ (.A(_21874_),
    .B(_21877_),
    .S(_03224_),
    .Z(_03317_));
 MUX2_X1 _26610_ (.A(_00553_),
    .B(_00549_),
    .S(_03224_),
    .Z(_03318_));
 MUX2_X1 _26611_ (.A(_03317_),
    .B(_03318_),
    .S(_03228_),
    .Z(_03319_));
 MUX2_X1 _26612_ (.A(_03282_),
    .B(_03286_),
    .S(_03274_),
    .Z(_03320_));
 MUX2_X1 _26613_ (.A(_03319_),
    .B(_03320_),
    .S(_03280_),
    .Z(_03321_));
 MUX2_X1 _26614_ (.A(_03316_),
    .B(_03321_),
    .S(_03299_),
    .Z(_03322_));
 AOI21_X2 _26615_ (.A(_03279_),
    .B1(_03302_),
    .B2(_03274_),
    .ZN(_03323_));
 NAND2_X1 _26616_ (.A1(_03299_),
    .A2(_03323_),
    .ZN(_03324_));
 MUX2_X1 _26617_ (.A(_03322_),
    .B(_03324_),
    .S(_03270_),
    .Z(_03325_));
 OR2_X1 _26618_ (.A1(_03309_),
    .A2(_03325_),
    .ZN(_14139_));
 INV_X1 _26619_ (.A(_14139_),
    .ZN(_14133_));
 NOR3_X4 _26620_ (.A1(_03198_),
    .A2(_03295_),
    .A3(_03296_),
    .ZN(_03326_));
 AOI21_X4 _26621_ (.A(_03197_),
    .B1(_03290_),
    .B2(_03292_),
    .ZN(_03327_));
 NOR2_X4 _26622_ (.A1(_03326_),
    .A2(_03327_),
    .ZN(_03328_));
 XNOR2_X2 _26623_ (.A(_03200_),
    .B(_03268_),
    .ZN(_03329_));
 NAND2_X1 _26624_ (.A1(_03257_),
    .A2(_03329_),
    .ZN(_03330_));
 NOR2_X1 _26625_ (.A1(_03328_),
    .A2(_03330_),
    .ZN(_03331_));
 NAND2_X1 _26626_ (.A1(_03323_),
    .A2(_03331_),
    .ZN(_21907_));
 INV_X1 _26627_ (.A(_21907_),
    .ZN(_21911_));
 OR3_X1 _26628_ (.A1(_03328_),
    .A2(_03304_),
    .A3(_03330_),
    .ZN(_21900_));
 INV_X1 _26629_ (.A(_21900_),
    .ZN(_21904_));
 MUX2_X1 _26630_ (.A(_21865_),
    .B(_21859_),
    .S(_03279_),
    .Z(_03332_));
 NOR2_X1 _26631_ (.A1(_03274_),
    .A2(_03279_),
    .ZN(_03333_));
 AOI22_X1 _26632_ (.A1(_03274_),
    .A2(_03332_),
    .B1(_03333_),
    .B2(_21862_),
    .ZN(_03334_));
 MUX2_X1 _26633_ (.A(_00554_),
    .B(_00557_),
    .S(_03279_),
    .Z(_03335_));
 AOI22_X1 _26634_ (.A1(_00558_),
    .A2(_03333_),
    .B1(_03335_),
    .B2(_03274_),
    .ZN(_03336_));
 MUX2_X1 _26635_ (.A(_03334_),
    .B(_03336_),
    .S(_03228_),
    .Z(_03337_));
 NAND2_X1 _26636_ (.A1(_03331_),
    .A2(_03337_),
    .ZN(_21935_));
 INV_X1 _26637_ (.A(_21935_),
    .ZN(_21939_));
 NAND2_X1 _26638_ (.A1(_03274_),
    .A2(_03280_),
    .ZN(_03338_));
 MUX2_X1 _26639_ (.A(_03275_),
    .B(_03303_),
    .S(_03279_),
    .Z(_03339_));
 MUX2_X1 _26640_ (.A(_03338_),
    .B(_03339_),
    .S(_03299_),
    .Z(_03340_));
 OR2_X1 _26641_ (.A1(_03330_),
    .A2(_03340_),
    .ZN(_21914_));
 INV_X1 _26642_ (.A(_21914_),
    .ZN(_21918_));
 NOR2_X1 _26643_ (.A1(_03309_),
    .A2(_03270_),
    .ZN(_03341_));
 NAND2_X1 _26644_ (.A1(_03328_),
    .A2(_03323_),
    .ZN(_03342_));
 OAI21_X1 _26645_ (.A(_03342_),
    .B1(_03316_),
    .B2(_03328_),
    .ZN(_03343_));
 AND2_X1 _26646_ (.A1(_03341_),
    .A2(_03343_),
    .ZN(_21921_));
 INV_X1 _26647_ (.A(_21921_),
    .ZN(_21925_));
 MUX2_X1 _26648_ (.A(_03281_),
    .B(_03304_),
    .S(_03328_),
    .Z(_03344_));
 NOR2_X1 _26649_ (.A1(_03330_),
    .A2(_03344_),
    .ZN(_21928_));
 INV_X1 _26650_ (.A(_21928_),
    .ZN(_21932_));
 NOR3_X1 _26651_ (.A1(_03280_),
    .A2(_03311_),
    .A3(_03313_),
    .ZN(_03345_));
 AOI21_X1 _26652_ (.A(_03345_),
    .B1(_03319_),
    .B2(_03280_),
    .ZN(_03346_));
 MUX2_X1 _26653_ (.A(_03337_),
    .B(_03346_),
    .S(_03299_),
    .Z(_03347_));
 AND2_X1 _26654_ (.A1(_03341_),
    .A2(_03347_),
    .ZN(_21945_));
 INV_X1 _26655_ (.A(_21945_),
    .ZN(_21949_));
 MUX2_X1 _26656_ (.A(_03284_),
    .B(_03285_),
    .S(_03329_),
    .Z(_03348_));
 NOR2_X1 _26657_ (.A1(_03279_),
    .A2(_03348_),
    .ZN(_03349_));
 NOR3_X1 _26658_ (.A1(_03280_),
    .A2(_03270_),
    .A3(_03278_),
    .ZN(_03350_));
 OAI21_X1 _26659_ (.A(_03299_),
    .B1(_03349_),
    .B2(_03350_),
    .ZN(_03351_));
 OR2_X1 _26660_ (.A1(_03270_),
    .A2(_03339_),
    .ZN(_03352_));
 OAI21_X1 _26661_ (.A(_03351_),
    .B1(_03352_),
    .B2(_03299_),
    .ZN(_03353_));
 NAND2_X1 _26662_ (.A1(_03257_),
    .A2(_03353_),
    .ZN(_21942_));
 INV_X1 _26663_ (.A(_21942_),
    .ZN(_21896_));
 INV_X1 _26664_ (.A(\g_reduce0[8].adder.a[15] ),
    .ZN(_03354_));
 NOR2_X1 _26665_ (.A1(_03354_),
    .A2(\g_reduce0[8].adder.b[15] ),
    .ZN(_03355_));
 AND2_X1 _26666_ (.A1(_03354_),
    .A2(\g_reduce0[8].adder.b[15] ),
    .ZN(_03356_));
 OR2_X1 _26667_ (.A1(_03355_),
    .A2(_03356_),
    .ZN(_03357_));
 CLKBUF_X3 _26668_ (.A(_03357_),
    .Z(_03358_));
 BUF_X4 _26669_ (.A(_03358_),
    .Z(_03359_));
 BUF_X2 _26670_ (.A(_21910_),
    .Z(_03360_));
 NOR2_X1 _26671_ (.A1(_21940_),
    .A2(_21905_),
    .ZN(_03361_));
 BUF_X2 _26672_ (.A(_21938_),
    .Z(_03362_));
 INV_X1 _26673_ (.A(_03362_),
    .ZN(_03363_));
 INV_X1 _26674_ (.A(_21898_),
    .ZN(_03364_));
 INV_X1 _26675_ (.A(_21899_),
    .ZN(_03365_));
 AOI21_X1 _26676_ (.A(_21892_),
    .B1(_14135_),
    .B2(_21893_),
    .ZN(_03366_));
 OAI21_X2 _26677_ (.A(_03364_),
    .B1(_03365_),
    .B2(_03366_),
    .ZN(_03367_));
 AND2_X1 _26678_ (.A1(_21948_),
    .A2(_03367_),
    .ZN(_03368_));
 INV_X1 _26679_ (.A(_21919_),
    .ZN(_03369_));
 INV_X1 _26680_ (.A(_21923_),
    .ZN(_03370_));
 NOR2_X1 _26681_ (.A1(_21930_),
    .A2(_21947_),
    .ZN(_03371_));
 NAND3_X1 _26682_ (.A1(_03369_),
    .A2(_03370_),
    .A3(_03371_),
    .ZN(_03372_));
 CLKBUF_X3 _26683_ (.A(_21917_),
    .Z(_03373_));
 CLKBUF_X3 _26684_ (.A(_21924_),
    .Z(_03374_));
 OAI21_X2 _26685_ (.A(_03374_),
    .B1(_21931_),
    .B2(_21930_),
    .ZN(_03375_));
 AOI21_X2 _26686_ (.A(_03373_),
    .B1(_03370_),
    .B2(_03375_),
    .ZN(_03376_));
 OAI221_X2 _26687_ (.A(_03363_),
    .B1(_03368_),
    .B2(_03372_),
    .C1(_03376_),
    .C2(_21919_),
    .ZN(_03377_));
 INV_X1 _26688_ (.A(_21905_),
    .ZN(_03378_));
 CLKBUF_X3 _26689_ (.A(_21903_),
    .Z(_03379_));
 AOI221_X2 _26690_ (.A(_03360_),
    .B1(_03361_),
    .B2(_03377_),
    .C1(_03378_),
    .C2(_03379_),
    .ZN(_03380_));
 NOR2_X2 _26691_ (.A1(_21912_),
    .A2(_03380_),
    .ZN(_03381_));
 NOR2_X1 _26692_ (.A1(_03359_),
    .A2(_03381_),
    .ZN(_03382_));
 NOR2_X2 _26693_ (.A1(_03284_),
    .A2(_03279_),
    .ZN(_03383_));
 NAND2_X4 _26694_ (.A1(_03298_),
    .A2(_03383_),
    .ZN(_03384_));
 NOR3_X4 _26695_ (.A1(_03309_),
    .A2(_03269_),
    .A3(_03384_),
    .ZN(_03385_));
 BUF_X1 _26696_ (.A(_21916_),
    .Z(_03386_));
 NOR2_X1 _26697_ (.A1(_03373_),
    .A2(_03386_),
    .ZN(_03387_));
 NOR2_X1 _26698_ (.A1(_21926_),
    .A2(_03386_),
    .ZN(_03388_));
 AOI21_X2 _26699_ (.A(_03387_),
    .B1(_03388_),
    .B2(_03374_),
    .ZN(_03389_));
 NOR3_X1 _26700_ (.A1(_21926_),
    .A2(_03386_),
    .A3(_21933_),
    .ZN(_03390_));
 INV_X1 _26701_ (.A(_21943_),
    .ZN(_03391_));
 INV_X1 _26702_ (.A(_21944_),
    .ZN(_03392_));
 AOI21_X1 _26703_ (.A(_21894_),
    .B1(_14138_),
    .B2(_21895_),
    .ZN(_03393_));
 OAI21_X1 _26704_ (.A(_03391_),
    .B1(_03392_),
    .B2(_03393_),
    .ZN(_03394_));
 INV_X1 _26705_ (.A(_21948_),
    .ZN(_03395_));
 AOI21_X1 _26706_ (.A(_21950_),
    .B1(_03394_),
    .B2(_03395_),
    .ZN(_03396_));
 OAI21_X2 _26707_ (.A(_03390_),
    .B1(_03396_),
    .B2(_21931_),
    .ZN(_03397_));
 AND3_X1 _26708_ (.A1(_03362_),
    .A2(_03389_),
    .A3(_03397_),
    .ZN(_03398_));
 BUF_X1 _26709_ (.A(_21902_),
    .Z(_03399_));
 OR3_X1 _26710_ (.A1(_21909_),
    .A2(_21937_),
    .A3(_03399_),
    .ZN(_03400_));
 OAI21_X1 _26711_ (.A(_03360_),
    .B1(_03399_),
    .B2(_03379_),
    .ZN(_03401_));
 INV_X1 _26712_ (.A(_03401_),
    .ZN(_03402_));
 OAI221_X2 _26713_ (.A(_03359_),
    .B1(_03398_),
    .B2(_03400_),
    .C1(_03402_),
    .C2(_21909_),
    .ZN(_03403_));
 AOI21_X4 _26714_ (.A(_03382_),
    .B1(_03385_),
    .B2(_03403_),
    .ZN(_03404_));
 XNOR2_X2 _26715_ (.A(\g_reduce0[8].adder.a[15] ),
    .B(\g_reduce0[8].adder.b[15] ),
    .ZN(_03405_));
 BUF_X4 _26716_ (.A(_03405_),
    .Z(_03406_));
 BUF_X4 _26717_ (.A(_03406_),
    .Z(_03407_));
 NOR2_X1 _26718_ (.A1(_21909_),
    .A2(_03407_),
    .ZN(_03408_));
 NOR3_X1 _26719_ (.A1(_03373_),
    .A2(_03362_),
    .A3(_03370_),
    .ZN(_03409_));
 NOR3_X1 _26720_ (.A1(_03373_),
    .A2(_03362_),
    .A3(_03375_),
    .ZN(_03410_));
 AOI21_X1 _26721_ (.A(_21898_),
    .B1(_14136_),
    .B2(_21899_),
    .ZN(_03411_));
 OAI21_X1 _26722_ (.A(_03371_),
    .B1(_03411_),
    .B2(_03395_),
    .ZN(_03412_));
 AOI221_X2 _26723_ (.A(_03409_),
    .B1(_03410_),
    .B2(_03412_),
    .C1(_21919_),
    .C2(_03363_),
    .ZN(_03413_));
 AOI22_X1 _26724_ (.A1(_03379_),
    .A2(_03378_),
    .B1(_03361_),
    .B2(_03413_),
    .ZN(_03414_));
 AOI21_X1 _26725_ (.A(_03408_),
    .B1(_03414_),
    .B2(_03407_),
    .ZN(_03415_));
 NOR3_X1 _26726_ (.A1(_21937_),
    .A2(_21926_),
    .A3(_03386_),
    .ZN(_03416_));
 INV_X1 _26727_ (.A(_21950_),
    .ZN(_03417_));
 AOI21_X1 _26728_ (.A(_21943_),
    .B1(_14140_),
    .B2(_21944_),
    .ZN(_03418_));
 OAI21_X1 _26729_ (.A(_03417_),
    .B1(_03418_),
    .B2(_21948_),
    .ZN(_03419_));
 INV_X1 _26730_ (.A(_21931_),
    .ZN(_03420_));
 AOI21_X2 _26731_ (.A(_21933_),
    .B1(_03419_),
    .B2(_03420_),
    .ZN(_03421_));
 OAI21_X2 _26732_ (.A(_03416_),
    .B1(_03421_),
    .B2(_03374_),
    .ZN(_03422_));
 OAI21_X1 _26733_ (.A(_03362_),
    .B1(_03386_),
    .B2(_03373_),
    .ZN(_03423_));
 INV_X1 _26734_ (.A(_21937_),
    .ZN(_03424_));
 AOI21_X2 _26735_ (.A(_03406_),
    .B1(_03423_),
    .B2(_03424_),
    .ZN(_03425_));
 AND3_X1 _26736_ (.A1(_03379_),
    .A2(_03422_),
    .A3(_03425_),
    .ZN(_03426_));
 NOR3_X1 _26737_ (.A1(_21909_),
    .A2(_03399_),
    .A3(_03407_),
    .ZN(_03427_));
 AOI21_X1 _26738_ (.A(_03427_),
    .B1(_03407_),
    .B2(_21912_),
    .ZN(_03428_));
 OAI22_X1 _26739_ (.A1(_03360_),
    .A2(_03415_),
    .B1(_03426_),
    .B2(_03428_),
    .ZN(_03429_));
 CLKBUF_X3 _26740_ (.A(_03429_),
    .Z(_03430_));
 INV_X2 _26741_ (.A(_03430_),
    .ZN(_03431_));
 XNOR2_X2 _26742_ (.A(_03385_),
    .B(_03431_),
    .ZN(_03432_));
 INV_X1 _26743_ (.A(_03399_),
    .ZN(_03433_));
 OAI21_X1 _26744_ (.A(_03424_),
    .B1(_03433_),
    .B2(_03405_),
    .ZN(_03434_));
 INV_X1 _26745_ (.A(_03379_),
    .ZN(_03435_));
 AOI21_X1 _26746_ (.A(_21905_),
    .B1(_03435_),
    .B2(_21940_),
    .ZN(_03436_));
 AOI221_X2 _26747_ (.A(_03434_),
    .B1(_03397_),
    .B2(_03389_),
    .C1(_03406_),
    .C2(_03436_),
    .ZN(_03437_));
 AND2_X1 _26748_ (.A1(_03405_),
    .A2(_03361_),
    .ZN(_03438_));
 NOR3_X1 _26749_ (.A1(_03362_),
    .A2(_21937_),
    .A3(_03405_),
    .ZN(_03439_));
 AOI21_X1 _26750_ (.A(_03439_),
    .B1(_03406_),
    .B2(_21905_),
    .ZN(_03440_));
 AOI221_X2 _26751_ (.A(_03438_),
    .B1(_03358_),
    .B2(_03399_),
    .C1(_03379_),
    .C2(_03440_),
    .ZN(_03441_));
 NOR3_X2 _26752_ (.A1(_03379_),
    .A2(_03358_),
    .A3(_03377_),
    .ZN(_03442_));
 NOR3_X4 _26753_ (.A1(_03437_),
    .A2(_03441_),
    .A3(_03442_),
    .ZN(_03443_));
 XNOR2_X1 _26754_ (.A(_03360_),
    .B(_03443_),
    .ZN(_03444_));
 NOR2_X1 _26755_ (.A1(_21940_),
    .A2(_03358_),
    .ZN(_03445_));
 AOI22_X4 _26756_ (.A1(_03422_),
    .A2(_03425_),
    .B1(_03445_),
    .B2(_03413_),
    .ZN(_03446_));
 XNOR2_X2 _26757_ (.A(_03379_),
    .B(_03446_),
    .ZN(_03447_));
 AND4_X1 _26758_ (.A1(_03362_),
    .A2(_03359_),
    .A3(_03389_),
    .A4(_03397_),
    .ZN(_03448_));
 NAND2_X1 _26759_ (.A1(_03363_),
    .A2(_03358_),
    .ZN(_03449_));
 AOI21_X2 _26760_ (.A(_03449_),
    .B1(_03397_),
    .B2(_03389_),
    .ZN(_03450_));
 NOR2_X1 _26761_ (.A1(_03362_),
    .A2(_03358_),
    .ZN(_03451_));
 NOR2_X1 _26762_ (.A1(_03363_),
    .A2(_03358_),
    .ZN(_03452_));
 OAI22_X1 _26763_ (.A1(_21919_),
    .A2(_03376_),
    .B1(_03372_),
    .B2(_03368_),
    .ZN(_03453_));
 MUX2_X1 _26764_ (.A(_03451_),
    .B(_03452_),
    .S(_03453_),
    .Z(_03454_));
 NOR3_X4 _26765_ (.A1(_03448_),
    .A2(_03450_),
    .A3(_03454_),
    .ZN(_03455_));
 OR2_X1 _26766_ (.A1(_21931_),
    .A2(_03396_),
    .ZN(_03456_));
 NOR2_X2 _26767_ (.A1(_21933_),
    .A2(_03406_),
    .ZN(_03457_));
 INV_X1 _26768_ (.A(_21930_),
    .ZN(_03458_));
 AOI21_X1 _26769_ (.A(_21947_),
    .B1(_03367_),
    .B2(_21948_),
    .ZN(_03459_));
 OAI21_X2 _26770_ (.A(_03458_),
    .B1(_03459_),
    .B2(_03420_),
    .ZN(_03460_));
 AOI22_X4 _26771_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_03460_),
    .B2(_03406_),
    .ZN(_03461_));
 XNOR2_X2 _26772_ (.A(_03374_),
    .B(_03461_),
    .ZN(_03462_));
 NOR2_X1 _26773_ (.A1(_03395_),
    .A2(_03411_),
    .ZN(_03463_));
 NOR3_X1 _26774_ (.A1(_21930_),
    .A2(_21947_),
    .A3(_03463_),
    .ZN(_03464_));
 OAI21_X2 _26775_ (.A(_03370_),
    .B1(_03375_),
    .B2(_03464_),
    .ZN(_03465_));
 OR2_X1 _26776_ (.A1(_03374_),
    .A2(_03421_),
    .ZN(_03466_));
 NOR2_X1 _26777_ (.A1(_21926_),
    .A2(_03406_),
    .ZN(_03467_));
 AOI22_X4 _26778_ (.A1(_03407_),
    .A2(_03465_),
    .B1(_03466_),
    .B2(_03467_),
    .ZN(_03468_));
 XNOR2_X2 _26779_ (.A(_03373_),
    .B(_03468_),
    .ZN(_03469_));
 AOI21_X4 _26780_ (.A(_03455_),
    .B1(_03462_),
    .B2(_03469_),
    .ZN(_03470_));
 OAI21_X4 _26781_ (.A(_03444_),
    .B1(_03447_),
    .B2(_03470_),
    .ZN(_03471_));
 XOR2_X2 _26782_ (.A(_03373_),
    .B(_03468_),
    .Z(_03472_));
 NOR2_X1 _26783_ (.A1(_21947_),
    .A2(_03463_),
    .ZN(_03473_));
 MUX2_X1 _26784_ (.A(_03419_),
    .B(_03473_),
    .S(_03406_),
    .Z(_03474_));
 XNOR2_X2 _26785_ (.A(_03420_),
    .B(_03474_),
    .ZN(_03475_));
 INV_X2 _26786_ (.A(_03475_),
    .ZN(_03476_));
 NOR2_X1 _26787_ (.A1(_03406_),
    .A2(_03394_),
    .ZN(_03477_));
 AOI21_X2 _26788_ (.A(_03477_),
    .B1(_03367_),
    .B2(_03406_),
    .ZN(_03478_));
 XNOR2_X2 _26789_ (.A(_03395_),
    .B(_03478_),
    .ZN(_03479_));
 INV_X1 _26790_ (.A(_03479_),
    .ZN(_03480_));
 XNOR2_X1 _26791_ (.A(_14140_),
    .B(_21944_),
    .ZN(_03481_));
 NAND2_X2 _26792_ (.A1(_03358_),
    .A2(_03481_),
    .ZN(_03482_));
 XOR2_X2 _26793_ (.A(_14136_),
    .B(_21899_),
    .Z(_03483_));
 OAI21_X4 _26794_ (.A(_03482_),
    .B1(_03483_),
    .B2(_03359_),
    .ZN(_03484_));
 AND2_X1 _26795_ (.A1(_14137_),
    .A2(_03407_),
    .ZN(_03485_));
 AOI21_X2 _26796_ (.A(_03485_),
    .B1(_03359_),
    .B2(_14141_),
    .ZN(_03486_));
 AOI21_X2 _26797_ (.A(_03480_),
    .B1(_03484_),
    .B2(_03486_),
    .ZN(_03487_));
 NOR4_X2 _26798_ (.A1(_03447_),
    .A2(_03472_),
    .A3(_03476_),
    .A4(_03487_),
    .ZN(_03488_));
 NOR2_X1 _26799_ (.A1(_03471_),
    .A2(_03488_),
    .ZN(_03489_));
 NOR3_X4 _26800_ (.A1(_03447_),
    .A2(_03472_),
    .A3(_03476_),
    .ZN(_03490_));
 NOR3_X2 _26801_ (.A1(_21954_),
    .A2(_03359_),
    .A3(_03483_),
    .ZN(_03491_));
 NAND2_X1 _26802_ (.A1(_03490_),
    .A2(_03491_),
    .ZN(_03492_));
 NAND2_X1 _26803_ (.A1(_03489_),
    .A2(_03492_),
    .ZN(_03493_));
 NOR2_X2 _26804_ (.A1(_21956_),
    .A2(_03482_),
    .ZN(_03494_));
 NAND2_X1 _26805_ (.A1(_03490_),
    .A2(_03494_),
    .ZN(_03495_));
 NAND2_X1 _26806_ (.A1(_03489_),
    .A2(_03495_),
    .ZN(_03496_));
 NAND2_X1 _26807_ (.A1(_03224_),
    .A2(_03279_),
    .ZN(_03497_));
 MUX2_X1 _26808_ (.A(_00548_),
    .B(_21880_),
    .S(_21888_),
    .Z(_03498_));
 OAI22_X1 _26809_ (.A1(_21883_),
    .A2(_03497_),
    .B1(_03498_),
    .B2(_03224_),
    .ZN(_03499_));
 NOR3_X1 _26810_ (.A1(_03237_),
    .A2(_03239_),
    .A3(_03499_),
    .ZN(_03500_));
 MUX2_X1 _26811_ (.A(_00547_),
    .B(_00550_),
    .S(_21888_),
    .Z(_03501_));
 OAI22_X1 _26812_ (.A1(_00546_),
    .A2(_03497_),
    .B1(_03501_),
    .B2(_03274_),
    .ZN(_03502_));
 AOI21_X1 _26813_ (.A(_03502_),
    .B1(_03227_),
    .B2(_03204_),
    .ZN(_03503_));
 OAI22_X1 _26814_ (.A1(_03326_),
    .A2(_03327_),
    .B1(_03500_),
    .B2(_03503_),
    .ZN(_03504_));
 OAI221_X1 _26815_ (.A(_03504_),
    .B1(_03346_),
    .B2(_03298_),
    .C1(_03307_),
    .C2(_03308_),
    .ZN(_03505_));
 OAI221_X1 _26816_ (.A(_03337_),
    .B1(_03327_),
    .B2(_03326_),
    .C1(_03307_),
    .C2(_03308_),
    .ZN(_03506_));
 MUX2_X2 _26817_ (.A(_03505_),
    .B(_03506_),
    .S(_03269_),
    .Z(_03507_));
 MUX2_X2 _26818_ (.A(_03493_),
    .B(_03496_),
    .S(_03507_),
    .Z(_03508_));
 NAND2_X2 _26819_ (.A1(_03432_),
    .A2(_03508_),
    .ZN(_03509_));
 NAND2_X2 _26820_ (.A1(_03404_),
    .A2(_03509_),
    .ZN(_21958_));
 INV_X2 _26821_ (.A(_21958_),
    .ZN(_21960_));
 INV_X1 _26822_ (.A(_21963_),
    .ZN(_03510_));
 OR2_X1 _26823_ (.A1(_03403_),
    .A2(_03429_),
    .ZN(_03511_));
 NOR4_X4 _26824_ (.A1(_03309_),
    .A2(_03269_),
    .A3(_03384_),
    .A4(_03511_),
    .ZN(_03512_));
 OAI21_X2 _26825_ (.A(_03430_),
    .B1(_03381_),
    .B2(_03359_),
    .ZN(_03513_));
 INV_X2 _26826_ (.A(_03513_),
    .ZN(_03514_));
 OR3_X4 _26827_ (.A1(_03309_),
    .A2(_03269_),
    .A3(_03384_),
    .ZN(_03515_));
 AOI211_X2 _26828_ (.A(_03510_),
    .B(_03512_),
    .C1(_03514_),
    .C2(_03515_),
    .ZN(_03516_));
 XNOR2_X2 _26829_ (.A(_03435_),
    .B(_03446_),
    .ZN(_03517_));
 NAND2_X1 _26830_ (.A1(_03479_),
    .A2(_03484_),
    .ZN(_03518_));
 OR3_X2 _26831_ (.A1(_03462_),
    .A2(_03476_),
    .A3(_03518_),
    .ZN(_03519_));
 NOR2_X2 _26832_ (.A1(_03455_),
    .A2(_03472_),
    .ZN(_03520_));
 NAND4_X4 _26833_ (.A1(_03444_),
    .A2(_03517_),
    .A3(_03519_),
    .A4(_03520_),
    .ZN(_03521_));
 NOR2_X1 _26834_ (.A1(_21963_),
    .A2(_03513_),
    .ZN(_03522_));
 NAND2_X1 _26835_ (.A1(_03521_),
    .A2(_03522_),
    .ZN(_03523_));
 AOI21_X1 _26836_ (.A(_03523_),
    .B1(_03329_),
    .B2(_03257_),
    .ZN(_03524_));
 NOR2_X1 _26837_ (.A1(_21963_),
    .A2(_03511_),
    .ZN(_03525_));
 NAND4_X1 _26838_ (.A1(_03299_),
    .A2(_03383_),
    .A3(_03521_),
    .A4(_03525_),
    .ZN(_03526_));
 NOR3_X1 _26839_ (.A1(_03309_),
    .A2(_03270_),
    .A3(_03526_),
    .ZN(_03527_));
 OAI211_X2 _26840_ (.A(_03521_),
    .B(_03522_),
    .C1(_03328_),
    .C2(_03338_),
    .ZN(_03528_));
 OAI21_X1 _26841_ (.A(_03528_),
    .B1(_03521_),
    .B2(_03510_),
    .ZN(_03529_));
 OR3_X2 _26842_ (.A1(_03524_),
    .A2(_03527_),
    .A3(_03529_),
    .ZN(_03530_));
 NOR2_X2 _26843_ (.A1(_03516_),
    .A2(_03530_),
    .ZN(_03531_));
 INV_X4 _26844_ (.A(_03531_),
    .ZN(_21983_));
 CLKBUF_X3 _26845_ (.A(_21959_),
    .Z(_03532_));
 CLKBUF_X3 _26846_ (.A(_03532_),
    .Z(_03533_));
 AOI21_X4 _26847_ (.A(_03512_),
    .B1(_03514_),
    .B2(_03515_),
    .ZN(_03534_));
 BUF_X4 _26848_ (.A(_03534_),
    .Z(_03535_));
 INV_X1 _26849_ (.A(_21954_),
    .ZN(_03536_));
 NOR2_X1 _26850_ (.A1(_03536_),
    .A2(_03359_),
    .ZN(_03537_));
 AOI21_X4 _26851_ (.A(_03537_),
    .B1(_03359_),
    .B2(_21956_),
    .ZN(_03538_));
 NAND3_X1 _26852_ (.A1(_03533_),
    .A2(_03535_),
    .A3(_03538_),
    .ZN(_03539_));
 NOR2_X2 _26853_ (.A1(_03385_),
    .A2(_03513_),
    .ZN(_03540_));
 NOR2_X1 _26854_ (.A1(_03500_),
    .A2(_03503_),
    .ZN(_03541_));
 AOI21_X1 _26855_ (.A(_03541_),
    .B1(_03297_),
    .B2(_03293_),
    .ZN(_03542_));
 MUX2_X1 _26856_ (.A(_03314_),
    .B(_03319_),
    .S(_03280_),
    .Z(_03543_));
 AOI221_X1 _26857_ (.A(_03542_),
    .B1(_03543_),
    .B2(_03328_),
    .C1(_03253_),
    .C2(_03256_),
    .ZN(_03544_));
 OAI21_X1 _26858_ (.A(_03337_),
    .B1(_03327_),
    .B2(_03326_),
    .ZN(_03545_));
 AOI21_X1 _26859_ (.A(_03545_),
    .B1(_03256_),
    .B2(_03253_),
    .ZN(_03546_));
 MUX2_X2 _26860_ (.A(_03544_),
    .B(_03546_),
    .S(_03270_),
    .Z(_03547_));
 XNOR2_X2 _26861_ (.A(_03407_),
    .B(_03547_),
    .ZN(_03548_));
 NOR2_X1 _26862_ (.A1(_03532_),
    .A2(_03548_),
    .ZN(_03549_));
 XNOR2_X2 _26863_ (.A(_03515_),
    .B(_03431_),
    .ZN(_03550_));
 XOR2_X2 _26864_ (.A(_03360_),
    .B(_03443_),
    .Z(_03551_));
 OR3_X2 _26865_ (.A1(_03448_),
    .A2(_03450_),
    .A3(_03454_),
    .ZN(_03552_));
 NAND2_X1 _26866_ (.A1(_03552_),
    .A2(_03469_),
    .ZN(_03553_));
 NOR4_X4 _26867_ (.A1(_03551_),
    .A2(_03447_),
    .A3(_03519_),
    .A4(_03553_),
    .ZN(_03554_));
 INV_X2 _26868_ (.A(_03554_),
    .ZN(_03555_));
 OR2_X1 _26869_ (.A1(_21956_),
    .A2(_03482_),
    .ZN(_03556_));
 NOR2_X1 _26870_ (.A1(_03551_),
    .A2(_03447_),
    .ZN(_03557_));
 MUX2_X2 _26871_ (.A(_14141_),
    .B(_14137_),
    .S(_03407_),
    .Z(_03558_));
 AOI21_X1 _26872_ (.A(_03518_),
    .B1(_03538_),
    .B2(_03558_),
    .ZN(_03559_));
 NOR3_X1 _26873_ (.A1(_03462_),
    .A2(_03476_),
    .A3(_03559_),
    .ZN(_03560_));
 AND4_X1 _26874_ (.A1(_03487_),
    .A2(_03557_),
    .A3(_03520_),
    .A4(_03560_),
    .ZN(_03561_));
 NAND2_X1 _26875_ (.A1(_03556_),
    .A2(_03561_),
    .ZN(_03562_));
 NAND3_X1 _26876_ (.A1(_03536_),
    .A2(_03407_),
    .A3(_03484_),
    .ZN(_03563_));
 NAND2_X1 _26877_ (.A1(_03563_),
    .A2(_03561_),
    .ZN(_03564_));
 MUX2_X2 _26878_ (.A(_03562_),
    .B(_03564_),
    .S(_03547_),
    .Z(_03565_));
 OAI221_X2 _26879_ (.A(_03404_),
    .B1(_03550_),
    .B2(_03555_),
    .C1(_03565_),
    .C2(_03534_),
    .ZN(_03566_));
 BUF_X2 _26880_ (.A(_14143_),
    .Z(_03567_));
 OAI221_X2 _26881_ (.A(_03567_),
    .B1(_03512_),
    .B2(_03540_),
    .C1(_03548_),
    .C2(_03508_),
    .ZN(_03568_));
 CLKBUF_X3 _26882_ (.A(_03531_),
    .Z(_03569_));
 OAI33_X1 _26883_ (.A1(_03512_),
    .A2(_03540_),
    .A3(_03549_),
    .B1(_03566_),
    .B2(_03568_),
    .B3(_03569_),
    .ZN(_03570_));
 AND2_X1 _26884_ (.A1(_03539_),
    .A2(_03570_),
    .ZN(_03571_));
 NAND3_X1 _26885_ (.A1(_03533_),
    .A2(_03558_),
    .A3(_03535_),
    .ZN(_03572_));
 MUX2_X2 _26886_ (.A(_21956_),
    .B(_21954_),
    .S(_03407_),
    .Z(_03573_));
 OAI21_X1 _26887_ (.A(_03535_),
    .B1(_03573_),
    .B2(_03533_),
    .ZN(_03574_));
 INV_X2 _26888_ (.A(_03567_),
    .ZN(_03575_));
 AND2_X1 _26889_ (.A1(_03489_),
    .A2(_03492_),
    .ZN(_03576_));
 AND2_X1 _26890_ (.A1(_03489_),
    .A2(_03495_),
    .ZN(_03577_));
 MUX2_X2 _26891_ (.A(_03576_),
    .B(_03577_),
    .S(_03507_),
    .Z(_03578_));
 XNOR2_X2 _26892_ (.A(_03359_),
    .B(_03547_),
    .ZN(_03579_));
 NOR4_X4 _26893_ (.A1(_03575_),
    .A2(_03578_),
    .A3(_03534_),
    .A4(_03579_),
    .ZN(_03580_));
 NAND3_X1 _26894_ (.A1(_03298_),
    .A2(_03383_),
    .A3(_03403_),
    .ZN(_03581_));
 OAI33_X1 _26895_ (.A1(_03355_),
    .A2(_03356_),
    .A3(_03381_),
    .B1(_03581_),
    .B2(_03309_),
    .B3(_03269_),
    .ZN(_03582_));
 CLKBUF_X3 _26896_ (.A(_03582_),
    .Z(_03583_));
 AOI21_X2 _26897_ (.A(_03583_),
    .B1(_03538_),
    .B2(_03567_),
    .ZN(_03584_));
 AOI21_X4 _26898_ (.A(_03580_),
    .B1(_03584_),
    .B2(_03509_),
    .ZN(_03585_));
 NAND4_X1 _26899_ (.A1(_03487_),
    .A2(_03557_),
    .A3(_03520_),
    .A4(_03560_),
    .ZN(_03586_));
 NOR2_X1 _26900_ (.A1(_03494_),
    .A2(_03586_),
    .ZN(_03587_));
 NOR2_X1 _26901_ (.A1(_03491_),
    .A2(_03586_),
    .ZN(_03588_));
 MUX2_X1 _26902_ (.A(_03587_),
    .B(_03588_),
    .S(_03547_),
    .Z(_03589_));
 NOR3_X4 _26903_ (.A1(_03534_),
    .A2(_03554_),
    .A3(_03589_),
    .ZN(_03590_));
 NAND2_X2 _26904_ (.A1(_21983_),
    .A2(_03590_),
    .ZN(_03591_));
 OAI21_X2 _26905_ (.A(_03574_),
    .B1(_03585_),
    .B2(_03591_),
    .ZN(_03592_));
 AND3_X1 _26906_ (.A1(_03571_),
    .A2(_03572_),
    .A3(_03592_),
    .ZN(_21966_));
 NOR4_X4 _26907_ (.A1(_03185_),
    .A2(\g_reduce0[8].adder.a[12] ),
    .A3(\g_reduce0[8].adder.a[14] ),
    .A4(_03187_),
    .ZN(_03593_));
 NAND2_X1 _26908_ (.A1(\g_reduce0[8].adder.b[0] ),
    .A2(_03593_),
    .ZN(_03594_));
 NAND2_X4 _26909_ (.A1(_03189_),
    .A2(_03192_),
    .ZN(_03595_));
 OR4_X1 _26910_ (.A1(\g_reduce0[8].adder.b[11] ),
    .A2(\g_reduce0[8].adder.b[12] ),
    .A3(_03190_),
    .A4(_03191_),
    .ZN(_03596_));
 BUF_X2 _26911_ (.A(_03596_),
    .Z(_03597_));
 NAND2_X1 _26912_ (.A1(_03189_),
    .A2(_03597_),
    .ZN(_03598_));
 CLKBUF_X3 _26913_ (.A(_03598_),
    .Z(_03599_));
 INV_X1 _26914_ (.A(_21968_),
    .ZN(_03600_));
 INV_X1 _26915_ (.A(_21961_),
    .ZN(_03601_));
 NOR3_X1 _26916_ (.A1(_03601_),
    .A2(_03569_),
    .A3(_03566_),
    .ZN(_03602_));
 OAI21_X1 _26917_ (.A(_03571_),
    .B1(_03602_),
    .B2(_03535_),
    .ZN(_03603_));
 NAND2_X1 _26918_ (.A1(_03572_),
    .A2(_03592_),
    .ZN(_03604_));
 MUX2_X1 _26919_ (.A(_03571_),
    .B(_03603_),
    .S(_03604_),
    .Z(_03605_));
 CLKBUF_X3 _26920_ (.A(_03567_),
    .Z(_03606_));
 NOR2_X2 _26921_ (.A1(_03447_),
    .A2(_03470_),
    .ZN(_03607_));
 NOR2_X1 _26922_ (.A1(_03551_),
    .A2(_03607_),
    .ZN(_03608_));
 AOI21_X1 _26923_ (.A(_03550_),
    .B1(_03444_),
    .B2(_03447_),
    .ZN(_03609_));
 OAI33_X1 _26924_ (.A1(_03469_),
    .A2(_03608_),
    .A3(_03534_),
    .B1(_03609_),
    .B2(_03583_),
    .B3(_03552_),
    .ZN(_03610_));
 AND3_X1 _26925_ (.A1(_03606_),
    .A2(_03569_),
    .A3(_03610_),
    .ZN(_03611_));
 NOR2_X1 _26926_ (.A1(_03471_),
    .A2(_03490_),
    .ZN(_03612_));
 NOR2_X1 _26927_ (.A1(_03431_),
    .A2(_03612_),
    .ZN(_03613_));
 NOR2_X1 _26928_ (.A1(_03430_),
    .A2(_03612_),
    .ZN(_03614_));
 MUX2_X1 _26929_ (.A(_03613_),
    .B(_03614_),
    .S(_03385_),
    .Z(_03615_));
 NOR2_X1 _26930_ (.A1(_03486_),
    .A2(_03615_),
    .ZN(_03616_));
 NAND3_X1 _26931_ (.A1(_03444_),
    .A2(_03479_),
    .A3(_03558_),
    .ZN(_03617_));
 MUX2_X1 _26932_ (.A(_03491_),
    .B(_03494_),
    .S(_03507_),
    .Z(_03618_));
 OAI33_X1 _26933_ (.A1(_03550_),
    .A2(_03578_),
    .A3(_03573_),
    .B1(_03617_),
    .B2(_03618_),
    .B3(_03607_),
    .ZN(_03619_));
 OAI21_X2 _26934_ (.A(_03575_),
    .B1(_03516_),
    .B2(_03530_),
    .ZN(_03620_));
 OAI21_X2 _26935_ (.A(_03579_),
    .B1(_03578_),
    .B2(_03550_),
    .ZN(_03621_));
 NOR2_X1 _26936_ (.A1(_21983_),
    .A2(_03621_),
    .ZN(_03622_));
 AOI21_X1 _26937_ (.A(_03471_),
    .B1(_03490_),
    .B2(_03491_),
    .ZN(_03623_));
 AOI21_X1 _26938_ (.A(_03471_),
    .B1(_03490_),
    .B2(_03494_),
    .ZN(_03624_));
 MUX2_X1 _26939_ (.A(_03623_),
    .B(_03624_),
    .S(_03507_),
    .Z(_03625_));
 OAI21_X2 _26940_ (.A(_03479_),
    .B1(_03625_),
    .B2(_03550_),
    .ZN(_03626_));
 OAI21_X1 _26941_ (.A(_03484_),
    .B1(_03615_),
    .B2(_03479_),
    .ZN(_03627_));
 AOI21_X1 _26942_ (.A(_03569_),
    .B1(_03626_),
    .B2(_03627_),
    .ZN(_03628_));
 CLKBUF_X3 _26943_ (.A(_03575_),
    .Z(_03629_));
 OAI33_X1 _26944_ (.A1(_03616_),
    .A2(_03619_),
    .A3(_03620_),
    .B1(_03622_),
    .B2(_03628_),
    .B3(_03629_),
    .ZN(_03630_));
 INV_X1 _26945_ (.A(_03566_),
    .ZN(_21987_));
 NOR2_X1 _26946_ (.A1(_03583_),
    .A2(_21987_),
    .ZN(_03631_));
 NAND2_X1 _26947_ (.A1(_03430_),
    .A2(_03551_),
    .ZN(_03632_));
 NAND2_X1 _26948_ (.A1(_03431_),
    .A2(_03551_),
    .ZN(_03633_));
 MUX2_X2 _26949_ (.A(_03632_),
    .B(_03633_),
    .S(_03385_),
    .Z(_03634_));
 OR2_X1 _26950_ (.A1(_03583_),
    .A2(_03475_),
    .ZN(_03635_));
 XOR2_X1 _26951_ (.A(_03374_),
    .B(_03461_),
    .Z(_03636_));
 OR2_X1 _26952_ (.A1(_03583_),
    .A2(_03636_),
    .ZN(_03637_));
 NOR2_X1 _26953_ (.A1(_03431_),
    .A2(_03489_),
    .ZN(_03638_));
 NOR2_X1 _26954_ (.A1(_03430_),
    .A2(_03489_),
    .ZN(_03639_));
 MUX2_X1 _26955_ (.A(_03638_),
    .B(_03639_),
    .S(_03385_),
    .Z(_03640_));
 NAND2_X1 _26956_ (.A1(_03607_),
    .A2(_03476_),
    .ZN(_03641_));
 OAI222_X2 _26957_ (.A1(_03634_),
    .A2(_03635_),
    .B1(_03637_),
    .B2(_03640_),
    .C1(_03641_),
    .C2(_03534_),
    .ZN(_03642_));
 OAI21_X1 _26958_ (.A(_03404_),
    .B1(_03550_),
    .B2(_03447_),
    .ZN(_03643_));
 NOR2_X1 _26959_ (.A1(_03444_),
    .A2(_03643_),
    .ZN(_03644_));
 MUX2_X1 _26960_ (.A(_03642_),
    .B(_03644_),
    .S(_21983_),
    .Z(_03645_));
 AOI221_X2 _26961_ (.A(_03611_),
    .B1(_03630_),
    .B2(_03631_),
    .C1(_03629_),
    .C2(_03645_),
    .ZN(_03646_));
 OAI22_X4 _26962_ (.A1(_03533_),
    .A2(_03404_),
    .B1(_03535_),
    .B2(_03646_),
    .ZN(_03647_));
 NOR2_X1 _26963_ (.A1(_03606_),
    .A2(_03621_),
    .ZN(_03648_));
 NAND3_X1 _26964_ (.A1(_03432_),
    .A2(_03508_),
    .A3(_03538_),
    .ZN(_03649_));
 OAI21_X1 _26965_ (.A(_03430_),
    .B1(_03471_),
    .B2(_03490_),
    .ZN(_03650_));
 OAI21_X1 _26966_ (.A(_03431_),
    .B1(_03471_),
    .B2(_03490_),
    .ZN(_03651_));
 MUX2_X1 _26967_ (.A(_03650_),
    .B(_03651_),
    .S(_03385_),
    .Z(_03652_));
 NOR2_X1 _26968_ (.A1(_03607_),
    .A2(_03617_),
    .ZN(_03653_));
 MUX2_X1 _26969_ (.A(_03563_),
    .B(_03556_),
    .S(_03507_),
    .Z(_03654_));
 AOI22_X1 _26970_ (.A1(_03558_),
    .A2(_03652_),
    .B1(_03653_),
    .B2(_03654_),
    .ZN(_03655_));
 AOI21_X1 _26971_ (.A(_03575_),
    .B1(_03649_),
    .B2(_03655_),
    .ZN(_03656_));
 NAND2_X2 _26972_ (.A1(_03569_),
    .A2(_03590_),
    .ZN(_03657_));
 NOR3_X1 _26973_ (.A1(_03648_),
    .A2(_03656_),
    .A3(_03657_),
    .ZN(_03658_));
 MUX2_X1 _26974_ (.A(_03462_),
    .B(_03472_),
    .S(_03532_),
    .Z(_03659_));
 NOR2_X1 _26975_ (.A1(_03403_),
    .A2(_03430_),
    .ZN(_03660_));
 MUX2_X2 _26976_ (.A(_03660_),
    .B(_03514_),
    .S(_03515_),
    .Z(_03661_));
 AND4_X2 _26977_ (.A1(_03661_),
    .A2(_03555_),
    .A3(_03530_),
    .A4(_03565_),
    .ZN(_03662_));
 NAND2_X1 _26978_ (.A1(_03606_),
    .A2(_03642_),
    .ZN(_03663_));
 NAND2_X1 _26979_ (.A1(_03629_),
    .A2(_03404_),
    .ZN(_03664_));
 NAND2_X1 _26980_ (.A1(_03626_),
    .A2(_03627_),
    .ZN(_03665_));
 OAI21_X2 _26981_ (.A(_03663_),
    .B1(_03664_),
    .B2(_03665_),
    .ZN(_03666_));
 AOI221_X2 _26982_ (.A(_03658_),
    .B1(_03659_),
    .B2(_03535_),
    .C1(_03662_),
    .C2(_03666_),
    .ZN(_03667_));
 NAND3_X4 _26983_ (.A1(_03661_),
    .A2(_03555_),
    .A3(_03565_),
    .ZN(_03668_));
 OR4_X1 _26984_ (.A1(_03668_),
    .A2(_03616_),
    .A3(_03619_),
    .A4(_03620_),
    .ZN(_03669_));
 NAND4_X1 _26985_ (.A1(_03606_),
    .A2(_03569_),
    .A3(_03590_),
    .A4(_03621_),
    .ZN(_03670_));
 MUX2_X1 _26986_ (.A(_03480_),
    .B(_03476_),
    .S(_03532_),
    .Z(_03671_));
 NAND2_X1 _26987_ (.A1(_03535_),
    .A2(_03671_),
    .ZN(_03672_));
 NAND4_X1 _26988_ (.A1(_03606_),
    .A2(_03662_),
    .A3(_03626_),
    .A4(_03627_),
    .ZN(_03673_));
 NAND4_X2 _26989_ (.A1(_03669_),
    .A2(_03670_),
    .A3(_03672_),
    .A4(_03673_),
    .ZN(_03674_));
 MUX2_X1 _26990_ (.A(_03476_),
    .B(_03462_),
    .S(_03532_),
    .Z(_03675_));
 OR3_X1 _26991_ (.A1(_03431_),
    .A2(_03479_),
    .A3(_03612_),
    .ZN(_03676_));
 OR3_X1 _26992_ (.A1(_03430_),
    .A2(_03479_),
    .A3(_03612_),
    .ZN(_03677_));
 MUX2_X1 _26993_ (.A(_03676_),
    .B(_03677_),
    .S(_03385_),
    .Z(_03678_));
 OAI221_X2 _26994_ (.A(_03430_),
    .B1(_03551_),
    .B2(_03607_),
    .C1(_03270_),
    .C2(_03309_),
    .ZN(_03679_));
 NOR3_X1 _26995_ (.A1(_03328_),
    .A2(_03338_),
    .A3(_03430_),
    .ZN(_03680_));
 NAND4_X1 _26996_ (.A1(_03257_),
    .A2(_03329_),
    .A3(_03471_),
    .A4(_03680_),
    .ZN(_03681_));
 AOI21_X1 _26997_ (.A(_03431_),
    .B1(_03383_),
    .B2(_03299_),
    .ZN(_03682_));
 AOI21_X1 _26998_ (.A(_03475_),
    .B1(_03682_),
    .B2(_03471_),
    .ZN(_03683_));
 NAND3_X2 _26999_ (.A1(_03679_),
    .A2(_03681_),
    .A3(_03683_),
    .ZN(_03684_));
 AOI211_X2 _27000_ (.A(_03575_),
    .B(_03583_),
    .C1(_03678_),
    .C2(_03684_),
    .ZN(_03685_));
 AOI22_X2 _27001_ (.A1(_03535_),
    .A2(_03675_),
    .B1(_03685_),
    .B2(_03662_),
    .ZN(_03686_));
 NOR2_X1 _27002_ (.A1(_03607_),
    .A2(_03488_),
    .ZN(_03687_));
 NAND2_X1 _27003_ (.A1(_03687_),
    .A2(_03492_),
    .ZN(_03688_));
 NAND2_X1 _27004_ (.A1(_03687_),
    .A2(_03495_),
    .ZN(_03689_));
 MUX2_X1 _27005_ (.A(_03688_),
    .B(_03689_),
    .S(_03507_),
    .Z(_03690_));
 AND3_X1 _27006_ (.A1(_03486_),
    .A2(_03661_),
    .A3(_03690_),
    .ZN(_03691_));
 OR2_X1 _27007_ (.A1(_03583_),
    .A2(_03558_),
    .ZN(_03692_));
 OAI33_X1 _27008_ (.A1(_03583_),
    .A2(_03484_),
    .A3(_03640_),
    .B1(_03692_),
    .B2(_03444_),
    .B3(_03550_),
    .ZN(_03693_));
 OAI21_X1 _27009_ (.A(_03662_),
    .B1(_03691_),
    .B2(_03693_),
    .ZN(_03694_));
 OAI221_X2 _27010_ (.A(_03686_),
    .B1(_03657_),
    .B2(_03585_),
    .C1(_03606_),
    .C2(_03694_),
    .ZN(_03695_));
 NAND2_X1 _27011_ (.A1(_03674_),
    .A2(_03695_),
    .ZN(_03696_));
 NOR2_X2 _27012_ (.A1(_03667_),
    .A2(_03696_),
    .ZN(_03697_));
 NAND2_X2 _27013_ (.A1(_21983_),
    .A2(_03566_),
    .ZN(_03698_));
 OR3_X1 _27014_ (.A1(_03551_),
    .A2(_03486_),
    .A3(_03690_),
    .ZN(_03699_));
 NAND3_X1 _27015_ (.A1(_03432_),
    .A2(_03538_),
    .A3(_03690_),
    .ZN(_03700_));
 AOI21_X1 _27016_ (.A(_03629_),
    .B1(_03699_),
    .B2(_03700_),
    .ZN(_03701_));
 OR4_X1 _27017_ (.A1(_03535_),
    .A2(_03648_),
    .A3(_03698_),
    .A4(_03701_),
    .ZN(_03702_));
 BUF_X4 _27018_ (.A(_03661_),
    .Z(_03703_));
 MUX2_X1 _27019_ (.A(_03444_),
    .B(_03432_),
    .S(_03532_),
    .Z(_03704_));
 NOR2_X1 _27020_ (.A1(_03703_),
    .A2(_03704_),
    .ZN(_03705_));
 NOR2_X1 _27021_ (.A1(_21983_),
    .A2(_03668_),
    .ZN(_03706_));
 MUX2_X1 _27022_ (.A(_03644_),
    .B(_03610_),
    .S(_03629_),
    .Z(_03707_));
 AOI221_X2 _27023_ (.A(_03705_),
    .B1(_03706_),
    .B2(_03666_),
    .C1(_03662_),
    .C2(_03707_),
    .ZN(_03708_));
 NAND2_X2 _27024_ (.A1(_03702_),
    .A2(_03708_),
    .ZN(_03709_));
 MUX2_X1 _27025_ (.A(_03469_),
    .B(_03552_),
    .S(_03532_),
    .Z(_03710_));
 NAND2_X1 _27026_ (.A1(_21961_),
    .A2(_03661_),
    .ZN(_03711_));
 OAI22_X4 _27027_ (.A1(_03661_),
    .A2(_03710_),
    .B1(_03698_),
    .B2(_03711_),
    .ZN(_03712_));
 AOI21_X1 _27028_ (.A(_03629_),
    .B1(_03569_),
    .B2(_03691_),
    .ZN(_03713_));
 OAI22_X2 _27029_ (.A1(_03558_),
    .A2(_03634_),
    .B1(_03640_),
    .B2(_03484_),
    .ZN(_03714_));
 NAND3_X1 _27030_ (.A1(_03404_),
    .A2(_03569_),
    .A3(_03714_),
    .ZN(_03715_));
 MUX2_X1 _27031_ (.A(_03636_),
    .B(_03469_),
    .S(_03509_),
    .Z(_03716_));
 OAI21_X1 _27032_ (.A(_03404_),
    .B1(_21983_),
    .B2(_03714_),
    .ZN(_03717_));
 OAI211_X2 _27033_ (.A(_03713_),
    .B(_03715_),
    .C1(_03716_),
    .C2(_03717_),
    .ZN(_03718_));
 NOR2_X1 _27034_ (.A1(_03567_),
    .A2(_03531_),
    .ZN(_03719_));
 NAND2_X1 _27035_ (.A1(_03678_),
    .A2(_03684_),
    .ZN(_03720_));
 NAND2_X1 _27036_ (.A1(_03404_),
    .A2(_03720_),
    .ZN(_03721_));
 NOR3_X2 _27037_ (.A1(_03578_),
    .A2(_03534_),
    .A3(_03579_),
    .ZN(_03722_));
 AOI21_X2 _27038_ (.A(_03722_),
    .B1(_03573_),
    .B2(_21960_),
    .ZN(_03723_));
 NOR2_X1 _27039_ (.A1(_03567_),
    .A2(_21983_),
    .ZN(_03724_));
 AOI221_X2 _27040_ (.A(_03668_),
    .B1(_03719_),
    .B2(_03721_),
    .C1(_03723_),
    .C2(_03724_),
    .ZN(_03725_));
 AOI21_X4 _27041_ (.A(_03712_),
    .B1(_03718_),
    .B2(_03725_),
    .ZN(_03726_));
 NAND3_X1 _27042_ (.A1(_03575_),
    .A2(_03569_),
    .A3(_03590_),
    .ZN(_03727_));
 NOR2_X1 _27043_ (.A1(_03691_),
    .A2(_03693_),
    .ZN(_03728_));
 MUX2_X1 _27044_ (.A(_03517_),
    .B(_03444_),
    .S(_21959_),
    .Z(_03729_));
 OAI222_X2 _27045_ (.A1(_03585_),
    .A2(_03698_),
    .B1(_03727_),
    .B2(_03728_),
    .C1(_03729_),
    .C2(_03661_),
    .ZN(_03730_));
 NOR2_X1 _27046_ (.A1(_03575_),
    .A2(_03668_),
    .ZN(_03731_));
 OR4_X1 _27047_ (.A1(_03309_),
    .A2(_03270_),
    .A3(_03384_),
    .A4(_03633_),
    .ZN(_03732_));
 OAI21_X1 _27048_ (.A(_03732_),
    .B1(_03632_),
    .B2(_03385_),
    .ZN(_03733_));
 OAI22_X1 _27049_ (.A1(_03550_),
    .A2(_03552_),
    .B1(_03733_),
    .B2(_03517_),
    .ZN(_03734_));
 MUX2_X1 _27050_ (.A(_03720_),
    .B(_03734_),
    .S(_21983_),
    .Z(_03735_));
 NOR2_X1 _27051_ (.A1(_03668_),
    .A2(_03620_),
    .ZN(_03736_));
 MUX2_X1 _27052_ (.A(_03462_),
    .B(_03472_),
    .S(_03509_),
    .Z(_03737_));
 AOI221_X2 _27053_ (.A(_03730_),
    .B1(_03731_),
    .B2(_03735_),
    .C1(_03736_),
    .C2(_03737_),
    .ZN(_03738_));
 NOR2_X1 _27054_ (.A1(_03629_),
    .A2(_03665_),
    .ZN(_03739_));
 NOR3_X1 _27055_ (.A1(_03606_),
    .A2(_03616_),
    .A3(_03619_),
    .ZN(_03740_));
 OAI21_X1 _27056_ (.A(_03706_),
    .B1(_03739_),
    .B2(_03740_),
    .ZN(_03741_));
 MUX2_X1 _27057_ (.A(_03552_),
    .B(_03517_),
    .S(_03532_),
    .Z(_03742_));
 OAI22_X2 _27058_ (.A1(_03568_),
    .A2(_03698_),
    .B1(_03742_),
    .B2(_03703_),
    .ZN(_03743_));
 MUX2_X1 _27059_ (.A(_03642_),
    .B(_03610_),
    .S(_03606_),
    .Z(_03744_));
 AOI21_X2 _27060_ (.A(_03743_),
    .B1(_03744_),
    .B2(_03662_),
    .ZN(_03745_));
 AOI211_X2 _27061_ (.A(_03726_),
    .B(_03738_),
    .C1(_03741_),
    .C2(_03745_),
    .ZN(_03746_));
 MUX2_X1 _27062_ (.A(_03484_),
    .B(_03479_),
    .S(_03532_),
    .Z(_03747_));
 OAI22_X2 _27063_ (.A1(_03601_),
    .A2(_03657_),
    .B1(_03747_),
    .B2(_03703_),
    .ZN(_03748_));
 NOR3_X1 _27064_ (.A1(_03629_),
    .A2(_03691_),
    .A3(_03693_),
    .ZN(_03749_));
 AOI211_X2 _27065_ (.A(_03591_),
    .B(_03749_),
    .C1(_03723_),
    .C2(_03629_),
    .ZN(_03750_));
 NOR2_X2 _27066_ (.A1(_03748_),
    .A2(_03750_),
    .ZN(_03751_));
 MUX2_X1 _27067_ (.A(_03558_),
    .B(_03484_),
    .S(_03532_),
    .Z(_03752_));
 OAI33_X1 _27068_ (.A1(_03591_),
    .A2(_03648_),
    .A3(_03656_),
    .B1(_03752_),
    .B2(_03512_),
    .B3(_03540_),
    .ZN(_21965_));
 NAND4_X2 _27069_ (.A1(_03571_),
    .A2(_03572_),
    .A3(_03592_),
    .A4(_21965_),
    .ZN(_03753_));
 NOR4_X1 _27070_ (.A1(_03629_),
    .A2(_03569_),
    .A3(_03668_),
    .A4(_03634_),
    .ZN(_03754_));
 NOR2_X1 _27071_ (.A1(_03606_),
    .A2(_03668_),
    .ZN(_03755_));
 AOI21_X1 _27072_ (.A(_03754_),
    .B1(_03755_),
    .B2(_03735_),
    .ZN(_03756_));
 MUX2_X1 _27073_ (.A(_03432_),
    .B(_03404_),
    .S(_03533_),
    .Z(_03757_));
 NAND3_X1 _27074_ (.A1(_03606_),
    .A2(_03706_),
    .A3(_03737_),
    .ZN(_03758_));
 AOI211_X2 _27075_ (.A(_03620_),
    .B(_03722_),
    .C1(_21960_),
    .C2(_03573_),
    .ZN(_03759_));
 OAI21_X1 _27076_ (.A(_03567_),
    .B1(_03516_),
    .B2(_03530_),
    .ZN(_03760_));
 OAI33_X1 _27077_ (.A1(_21961_),
    .A2(_03516_),
    .A3(_03530_),
    .B1(_03760_),
    .B2(_03691_),
    .B3(_03693_),
    .ZN(_03761_));
 OR4_X1 _27078_ (.A1(_03583_),
    .A2(_21987_),
    .A3(_03759_),
    .A4(_03761_),
    .ZN(_03762_));
 AND4_X1 _27079_ (.A1(_03756_),
    .A2(_03757_),
    .A3(_03758_),
    .A4(_03762_),
    .ZN(_03763_));
 NOR3_X1 _27080_ (.A1(_03751_),
    .A2(_03753_),
    .A3(_03763_),
    .ZN(_03764_));
 NAND4_X2 _27081_ (.A1(_03697_),
    .A2(_03709_),
    .A3(_03746_),
    .A4(_03764_),
    .ZN(_03765_));
 XOR2_X2 _27082_ (.A(_03647_),
    .B(_03765_),
    .Z(_03766_));
 MUX2_X1 _27083_ (.A(_03600_),
    .B(_03605_),
    .S(_03766_),
    .Z(_03767_));
 OAI221_X2 _27084_ (.A(_03594_),
    .B1(_03595_),
    .B2(_03212_),
    .C1(_03599_),
    .C2(_03767_),
    .ZN(_00112_));
 XNOR2_X1 _27085_ (.A(_21967_),
    .B(_03751_),
    .ZN(_03768_));
 NOR2_X1 _27086_ (.A1(_03598_),
    .A2(_03768_),
    .ZN(_03769_));
 NOR2_X1 _27087_ (.A1(_21968_),
    .A2(_03599_),
    .ZN(_03770_));
 MUX2_X1 _27088_ (.A(_03769_),
    .B(_03770_),
    .S(_03766_),
    .Z(_03771_));
 BUF_X4 _27089_ (.A(_03189_),
    .Z(_03772_));
 OAI22_X2 _27090_ (.A1(\g_reduce0[8].adder.b[1] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[1] ),
    .ZN(_03773_));
 NOR2_X1 _27091_ (.A1(_03771_),
    .A2(_03773_),
    .ZN(_00119_));
 OAI22_X2 _27092_ (.A1(\g_reduce0[8].adder.b[2] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[2] ),
    .ZN(_03774_));
 NOR2_X1 _27093_ (.A1(_03751_),
    .A2(_03753_),
    .ZN(_03775_));
 XOR2_X1 _27094_ (.A(_03674_),
    .B(_03775_),
    .Z(_03776_));
 NOR2_X1 _27095_ (.A1(_03599_),
    .A2(_03776_),
    .ZN(_03777_));
 INV_X4 _27096_ (.A(_03766_),
    .ZN(_21972_));
 MUX2_X1 _27097_ (.A(_03769_),
    .B(_03777_),
    .S(_21972_),
    .Z(_03778_));
 NOR2_X1 _27098_ (.A1(_03774_),
    .A2(_03778_),
    .ZN(_00120_));
 NOR2_X1 _27099_ (.A1(_03593_),
    .A2(_03192_),
    .ZN(_03779_));
 OR2_X1 _27100_ (.A1(_03748_),
    .A2(_03750_),
    .ZN(_03780_));
 NAND3_X1 _27101_ (.A1(_21967_),
    .A2(_03674_),
    .A3(_03780_),
    .ZN(_03781_));
 XOR2_X2 _27102_ (.A(_03695_),
    .B(_03781_),
    .Z(_03782_));
 AND2_X1 _27103_ (.A1(_03779_),
    .A2(_03782_),
    .ZN(_03783_));
 MUX2_X1 _27104_ (.A(_03777_),
    .B(_03783_),
    .S(_21972_),
    .Z(_03784_));
 OAI22_X2 _27105_ (.A1(\g_reduce0[8].adder.b[3] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[3] ),
    .ZN(_03785_));
 NOR2_X1 _27106_ (.A1(_03784_),
    .A2(_03785_),
    .ZN(_00121_));
 OAI22_X2 _27107_ (.A1(\g_reduce0[8].adder.b[4] ),
    .A2(_03189_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[4] ),
    .ZN(_03786_));
 NOR3_X1 _27108_ (.A1(_03696_),
    .A2(_03751_),
    .A3(_03753_),
    .ZN(_03787_));
 XOR2_X2 _27109_ (.A(_03667_),
    .B(_03787_),
    .Z(_03788_));
 OAI21_X1 _27110_ (.A(_03788_),
    .B1(_03782_),
    .B2(_03765_),
    .ZN(_03789_));
 NOR2_X1 _27111_ (.A1(_03647_),
    .A2(_03782_),
    .ZN(_03790_));
 AOI22_X1 _27112_ (.A1(_03647_),
    .A2(_03789_),
    .B1(_03790_),
    .B2(_03765_),
    .ZN(_03791_));
 AOI21_X1 _27113_ (.A(_03786_),
    .B1(_03791_),
    .B2(_03779_),
    .ZN(_00122_));
 OAI21_X1 _27114_ (.A(_03779_),
    .B1(_03647_),
    .B2(_03788_),
    .ZN(_03792_));
 INV_X1 _27115_ (.A(_21967_),
    .ZN(_03793_));
 NOR2_X1 _27116_ (.A1(_03793_),
    .A2(_03751_),
    .ZN(_03794_));
 NAND2_X1 _27117_ (.A1(_03697_),
    .A2(_03794_),
    .ZN(_03795_));
 XOR2_X2 _27118_ (.A(_03726_),
    .B(_03795_),
    .Z(_03796_));
 AOI21_X1 _27119_ (.A(_03792_),
    .B1(_03796_),
    .B2(_21972_),
    .ZN(_03797_));
 OAI22_X2 _27120_ (.A1(\g_reduce0[8].adder.b[5] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[5] ),
    .ZN(_03798_));
 NOR2_X1 _27121_ (.A1(_03797_),
    .A2(_03798_),
    .ZN(_00123_));
 NAND2_X1 _27122_ (.A1(_03741_),
    .A2(_03745_),
    .ZN(_03799_));
 NOR3_X1 _27123_ (.A1(_03667_),
    .A2(_03696_),
    .A3(_03726_),
    .ZN(_03800_));
 NAND2_X1 _27124_ (.A1(_03800_),
    .A2(_03775_),
    .ZN(_03801_));
 XNOR2_X1 _27125_ (.A(_03799_),
    .B(_03801_),
    .ZN(_03802_));
 NOR3_X1 _27126_ (.A1(_03599_),
    .A2(_03766_),
    .A3(_03802_),
    .ZN(_03803_));
 NOR3_X1 _27127_ (.A1(_03599_),
    .A2(_21972_),
    .A3(_03796_),
    .ZN(_03804_));
 OAI22_X2 _27128_ (.A1(\g_reduce0[8].adder.b[6] ),
    .A2(_03189_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[6] ),
    .ZN(_03805_));
 NOR3_X1 _27129_ (.A1(_03803_),
    .A2(_03804_),
    .A3(_03805_),
    .ZN(_00124_));
 OAI22_X2 _27130_ (.A1(\g_reduce0[8].adder.b[7] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[7] ),
    .ZN(_03806_));
 NOR3_X1 _27131_ (.A1(_03599_),
    .A2(_21972_),
    .A3(_03802_),
    .ZN(_03807_));
 NAND3_X1 _27132_ (.A1(_03800_),
    .A2(_03799_),
    .A3(_03794_),
    .ZN(_03808_));
 XOR2_X2 _27133_ (.A(_03738_),
    .B(_03808_),
    .Z(_03809_));
 NOR3_X1 _27134_ (.A1(_03599_),
    .A2(_03766_),
    .A3(_03809_),
    .ZN(_03810_));
 NOR3_X1 _27135_ (.A1(_03806_),
    .A2(_03807_),
    .A3(_03810_),
    .ZN(_00125_));
 OAI22_X2 _27136_ (.A1(\g_reduce0[8].adder.b[8] ),
    .A2(_03772_),
    .B1(_03595_),
    .B2(\g_reduce0[8].adder.a[8] ),
    .ZN(_03811_));
 NAND3_X1 _27137_ (.A1(_03697_),
    .A2(_03746_),
    .A3(_03775_),
    .ZN(_03812_));
 XNOR2_X1 _27138_ (.A(_03709_),
    .B(_03812_),
    .ZN(_03813_));
 NOR3_X1 _27139_ (.A1(_03599_),
    .A2(_03766_),
    .A3(_03813_),
    .ZN(_03814_));
 NOR3_X1 _27140_ (.A1(_03599_),
    .A2(_21972_),
    .A3(_03809_),
    .ZN(_03815_));
 NOR3_X1 _27141_ (.A1(_03811_),
    .A2(_03814_),
    .A3(_03815_),
    .ZN(_00126_));
 NOR2_X1 _27142_ (.A1(_03593_),
    .A2(_03597_),
    .ZN(_03816_));
 AOI22_X1 _27143_ (.A1(\g_reduce0[8].adder.b[9] ),
    .A2(_03593_),
    .B1(_03816_),
    .B2(\g_reduce0[8].adder.a[9] ),
    .ZN(_03817_));
 NAND3_X1 _27144_ (.A1(_03702_),
    .A2(_03708_),
    .A3(_03812_),
    .ZN(_03818_));
 NOR2_X1 _27145_ (.A1(_03599_),
    .A2(_03647_),
    .ZN(_03819_));
 OAI21_X1 _27146_ (.A(_03709_),
    .B1(_03763_),
    .B2(_03794_),
    .ZN(_03820_));
 OR2_X1 _27147_ (.A1(_03812_),
    .A2(_03820_),
    .ZN(_03821_));
 NAND3_X1 _27148_ (.A1(_03818_),
    .A2(_03819_),
    .A3(_03821_),
    .ZN(_03822_));
 AND2_X1 _27149_ (.A1(_03779_),
    .A2(_03647_),
    .ZN(_03823_));
 NAND4_X1 _27150_ (.A1(_03756_),
    .A2(_03757_),
    .A3(_03758_),
    .A4(_03762_),
    .ZN(_03824_));
 NOR3_X1 _27151_ (.A1(_03793_),
    .A2(_03751_),
    .A3(_03824_),
    .ZN(_03825_));
 AND4_X1 _27152_ (.A1(_03697_),
    .A2(_03709_),
    .A3(_03746_),
    .A4(_03825_),
    .ZN(_03826_));
 AOI21_X1 _27153_ (.A(_03751_),
    .B1(_03753_),
    .B2(_03793_),
    .ZN(_03827_));
 NAND4_X1 _27154_ (.A1(_03697_),
    .A2(_03709_),
    .A3(_03746_),
    .A4(_03827_),
    .ZN(_03828_));
 AND2_X1 _27155_ (.A1(_03824_),
    .A2(_03828_),
    .ZN(_03829_));
 OAI21_X1 _27156_ (.A(_03823_),
    .B1(_03826_),
    .B2(_03829_),
    .ZN(_03830_));
 NAND3_X1 _27157_ (.A1(_03817_),
    .A2(_03822_),
    .A3(_03830_),
    .ZN(_00127_));
 INV_X1 _27158_ (.A(_21975_),
    .ZN(_21969_));
 MUX2_X1 _27159_ (.A(_03186_),
    .B(_21974_),
    .S(_03597_),
    .Z(_03831_));
 MUX2_X1 _27160_ (.A(\g_reduce0[8].adder.b[10] ),
    .B(_03831_),
    .S(_03772_),
    .Z(_00113_));
 MUX2_X1 _27161_ (.A(_03185_),
    .B(_21982_),
    .S(_03597_),
    .Z(_03832_));
 MUX2_X1 _27162_ (.A(\g_reduce0[8].adder.b[11] ),
    .B(_03832_),
    .S(_03772_),
    .Z(_00114_));
 MUX2_X2 _27163_ (.A(_21850_),
    .B(_00556_),
    .S(_03240_),
    .Z(_03833_));
 NAND2_X1 _27164_ (.A1(_03533_),
    .A2(_21976_),
    .ZN(_03834_));
 XOR2_X1 _27165_ (.A(_03833_),
    .B(_03834_),
    .Z(_03835_));
 XOR2_X1 _27166_ (.A(_14145_),
    .B(_21986_),
    .Z(_03836_));
 MUX2_X1 _27167_ (.A(_03835_),
    .B(_03836_),
    .S(_03703_),
    .Z(_03837_));
 XOR2_X1 _27168_ (.A(_21981_),
    .B(_03837_),
    .Z(_03838_));
 MUX2_X1 _27169_ (.A(\g_reduce0[8].adder.a[12] ),
    .B(_03838_),
    .S(_03597_),
    .Z(_03839_));
 MUX2_X1 _27170_ (.A(\g_reduce0[8].adder.b[12] ),
    .B(_03839_),
    .S(_03772_),
    .Z(_00115_));
 INV_X1 _27171_ (.A(_14147_),
    .ZN(_14142_));
 MUX2_X1 _27172_ (.A(_21847_),
    .B(_00559_),
    .S(_03240_),
    .Z(_03840_));
 MUX2_X1 _27173_ (.A(_21853_),
    .B(_00551_),
    .S(_03240_),
    .Z(_03841_));
 NAND2_X1 _27174_ (.A1(_03533_),
    .A2(_21975_),
    .ZN(_03842_));
 NOR3_X1 _27175_ (.A1(_03833_),
    .A2(_03841_),
    .A3(_03842_),
    .ZN(_03843_));
 XNOR2_X1 _27176_ (.A(_03840_),
    .B(_03843_),
    .ZN(_03844_));
 INV_X1 _27177_ (.A(_21978_),
    .ZN(_03845_));
 INV_X1 _27178_ (.A(_21979_),
    .ZN(_03846_));
 OAI21_X1 _27179_ (.A(_03845_),
    .B1(_03846_),
    .B2(_14147_),
    .ZN(_03847_));
 AOI21_X1 _27180_ (.A(_21985_),
    .B1(_03847_),
    .B2(_21986_),
    .ZN(_03848_));
 XNOR2_X1 _27181_ (.A(_21990_),
    .B(_03848_),
    .ZN(_03849_));
 MUX2_X1 _27182_ (.A(_03844_),
    .B(_03849_),
    .S(_03703_),
    .Z(_03850_));
 NAND2_X1 _27183_ (.A1(_03533_),
    .A2(_21977_),
    .ZN(_03851_));
 OAI21_X1 _27184_ (.A(_03851_),
    .B1(_03841_),
    .B2(_03533_),
    .ZN(_03852_));
 MUX2_X1 _27185_ (.A(_14146_),
    .B(_03852_),
    .S(_03535_),
    .Z(_21980_));
 NAND3_X1 _27186_ (.A1(_21973_),
    .A2(_03837_),
    .A3(_21980_),
    .ZN(_03853_));
 XNOR2_X1 _27187_ (.A(_03850_),
    .B(_03853_),
    .ZN(_03854_));
 MUX2_X1 _27188_ (.A(\g_reduce0[8].adder.a[13] ),
    .B(_03854_),
    .S(_03597_),
    .Z(_03855_));
 MUX2_X1 _27189_ (.A(\g_reduce0[8].adder.b[13] ),
    .B(_03855_),
    .S(_03772_),
    .Z(_00116_));
 OR2_X1 _27190_ (.A1(_03190_),
    .A2(_03228_),
    .ZN(_03856_));
 NAND2_X1 _27191_ (.A1(\g_reduce0[8].adder.a[14] ),
    .A2(_03856_),
    .ZN(_03857_));
 NOR4_X1 _27192_ (.A1(_03703_),
    .A2(_03833_),
    .A3(_03834_),
    .A4(_03840_),
    .ZN(_03858_));
 AOI21_X1 _27193_ (.A(_21985_),
    .B1(_21986_),
    .B2(_14145_),
    .ZN(_03859_));
 INV_X1 _27194_ (.A(_03859_),
    .ZN(_03860_));
 AOI21_X1 _27195_ (.A(_21989_),
    .B1(_03860_),
    .B2(_21990_),
    .ZN(_03861_));
 AOI21_X1 _27196_ (.A(_03858_),
    .B1(_03861_),
    .B2(_03703_),
    .ZN(_03862_));
 NAND3_X1 _27197_ (.A1(_21981_),
    .A2(_03837_),
    .A3(_03850_),
    .ZN(_03863_));
 XOR2_X2 _27198_ (.A(_03862_),
    .B(_03863_),
    .Z(_03864_));
 MUX2_X1 _27199_ (.A(_03856_),
    .B(_03857_),
    .S(_03864_),
    .Z(_03865_));
 OAI22_X1 _27200_ (.A1(_03190_),
    .A2(_03189_),
    .B1(_03192_),
    .B2(_03865_),
    .ZN(_03866_));
 NOR2_X1 _27201_ (.A1(\g_reduce0[8].adder.a[14] ),
    .A2(_03593_),
    .ZN(_03867_));
 NAND3_X1 _27202_ (.A1(_03190_),
    .A2(_03272_),
    .A3(_03864_),
    .ZN(_03868_));
 OR2_X1 _27203_ (.A1(_03272_),
    .A2(_03864_),
    .ZN(_03869_));
 NAND3_X1 _27204_ (.A1(_03597_),
    .A2(_03868_),
    .A3(_03869_),
    .ZN(_03870_));
 AOI21_X1 _27205_ (.A(_03866_),
    .B1(_03867_),
    .B2(_03870_),
    .ZN(_00117_));
 OR2_X1 _27206_ (.A1(\g_reduce0[0].adder.x[10] ),
    .A2(\g_reduce0[0].adder.x[13] ),
    .ZN(_03871_));
 OR4_X1 _27207_ (.A1(\g_reduce0[0].adder.x[11] ),
    .A2(\g_reduce0[0].adder.x[12] ),
    .A3(\g_reduce0[0].adder.x[14] ),
    .A4(_03871_),
    .ZN(_03872_));
 CLKBUF_X3 _27208_ (.A(_03872_),
    .Z(_03873_));
 OR3_X1 _27209_ (.A1(\g_reduce0[2].adder.x[11] ),
    .A2(\g_reduce0[2].adder.x[10] ),
    .A3(\g_reduce0[2].adder.x[13] ),
    .ZN(_03874_));
 NOR3_X4 _27210_ (.A1(\g_reduce0[2].adder.x[12] ),
    .A2(\g_reduce0[2].adder.x[14] ),
    .A3(_03874_),
    .ZN(_03875_));
 CLKBUF_X3 _27211_ (.A(_22035_),
    .Z(_03876_));
 AOI21_X1 _27212_ (.A(_22034_),
    .B1(_21992_),
    .B2(_03876_),
    .ZN(_03877_));
 INV_X1 _27213_ (.A(_21998_),
    .ZN(_03878_));
 INV_X1 _27214_ (.A(_21999_),
    .ZN(_03879_));
 OAI21_X1 _27215_ (.A(_03878_),
    .B1(_22001_),
    .B2(_03879_),
    .ZN(_03880_));
 BUF_X4 _27216_ (.A(_21996_),
    .Z(_03881_));
 AOI21_X1 _27217_ (.A(_21995_),
    .B1(_03880_),
    .B2(_03881_),
    .ZN(_03882_));
 BUF_X4 _27218_ (.A(_21993_),
    .Z(_03883_));
 NAND2_X2 _27219_ (.A1(_22035_),
    .A2(_03883_),
    .ZN(_03884_));
 OAI21_X2 _27220_ (.A(_03877_),
    .B1(_03882_),
    .B2(_03884_),
    .ZN(_03885_));
 BUF_X2 _27221_ (.A(_22002_),
    .Z(_03886_));
 INV_X2 _27222_ (.A(_03886_),
    .ZN(_03887_));
 NAND2_X1 _27223_ (.A1(_03881_),
    .A2(_21999_),
    .ZN(_03888_));
 OR4_X1 _27224_ (.A1(_22004_),
    .A2(_03887_),
    .A3(_03888_),
    .A4(_03884_),
    .ZN(_03889_));
 INV_X1 _27225_ (.A(_22007_),
    .ZN(_03890_));
 AOI21_X1 _27226_ (.A(_22010_),
    .B1(_22011_),
    .B2(_22013_),
    .ZN(_03891_));
 INV_X1 _27227_ (.A(_22008_),
    .ZN(_03892_));
 OAI21_X2 _27228_ (.A(_03890_),
    .B1(_03891_),
    .B2(_03892_),
    .ZN(_03893_));
 AOI21_X1 _27229_ (.A(_03889_),
    .B1(_03893_),
    .B2(_22005_),
    .ZN(_03894_));
 INV_X1 _27230_ (.A(_03894_),
    .ZN(_03895_));
 NAND4_X2 _27231_ (.A1(_22005_),
    .A2(_22008_),
    .A3(_22011_),
    .A4(_22014_),
    .ZN(_03896_));
 AND3_X1 _27232_ (.A1(_22017_),
    .A2(_22020_),
    .A3(_22023_),
    .ZN(_03897_));
 INV_X1 _27233_ (.A(_22029_),
    .ZN(_03898_));
 INV_X1 _27234_ (.A(\g_reduce0[2].adder.x[0] ),
    .ZN(_03899_));
 AOI21_X1 _27235_ (.A(_03898_),
    .B1(_03899_),
    .B2(\g_reduce0[0].adder.x[0] ),
    .ZN(_03900_));
 OR2_X1 _27236_ (.A1(_22025_),
    .A2(_22028_),
    .ZN(_03901_));
 OAI221_X2 _27237_ (.A(_03897_),
    .B1(_03900_),
    .B2(_03901_),
    .C1(_22026_),
    .C2(_22025_),
    .ZN(_03902_));
 AOI21_X1 _27238_ (.A(_22019_),
    .B1(_22022_),
    .B2(_22020_),
    .ZN(_03903_));
 INV_X1 _27239_ (.A(_03903_),
    .ZN(_03904_));
 AOI21_X2 _27240_ (.A(_22016_),
    .B1(_03904_),
    .B2(_22017_),
    .ZN(_03905_));
 AOI21_X4 _27241_ (.A(_03896_),
    .B1(_03902_),
    .B2(_03905_),
    .ZN(_03906_));
 OAI21_X1 _27242_ (.A(_03885_),
    .B1(_03895_),
    .B2(_03906_),
    .ZN(_03907_));
 BUF_X4 _27243_ (.A(_03907_),
    .Z(_03908_));
 OAI21_X1 _27244_ (.A(_03873_),
    .B1(_03875_),
    .B2(_03908_),
    .ZN(_03909_));
 MUX2_X1 _27245_ (.A(\g_reduce0[0].adder.x[15] ),
    .B(\g_reduce0[2].adder.x[15] ),
    .S(_03909_),
    .Z(_00134_));
 INV_X2 _27246_ (.A(_03876_),
    .ZN(_03910_));
 INV_X2 _27247_ (.A(_03883_),
    .ZN(_03911_));
 NOR2_X2 _27248_ (.A1(_03910_),
    .A2(_03911_),
    .ZN(_03912_));
 INV_X1 _27249_ (.A(_21995_),
    .ZN(_03913_));
 INV_X1 _27250_ (.A(_22001_),
    .ZN(_03914_));
 AOI21_X1 _27251_ (.A(_21998_),
    .B1(_03914_),
    .B2(_21999_),
    .ZN(_03915_));
 INV_X2 _27252_ (.A(_21996_),
    .ZN(_03916_));
 OAI21_X1 _27253_ (.A(_03913_),
    .B1(_03915_),
    .B2(_03916_),
    .ZN(_03917_));
 AOI221_X2 _27254_ (.A(_22034_),
    .B1(_03912_),
    .B2(_03917_),
    .C1(_21992_),
    .C2(_03876_),
    .ZN(_03918_));
 AND4_X1 _27255_ (.A1(_22005_),
    .A2(_22008_),
    .A3(_22011_),
    .A4(_22014_),
    .ZN(_03919_));
 OAI21_X1 _27256_ (.A(_03897_),
    .B1(_22026_),
    .B2(_22025_),
    .ZN(_03920_));
 NOR2_X1 _27257_ (.A1(_22025_),
    .A2(_22028_),
    .ZN(_03921_));
 INV_X1 _27258_ (.A(\g_reduce0[0].adder.x[0] ),
    .ZN(_03922_));
 OAI21_X1 _27259_ (.A(_22029_),
    .B1(\g_reduce0[2].adder.x[0] ),
    .B2(_03922_),
    .ZN(_03923_));
 AOI21_X1 _27260_ (.A(_03920_),
    .B1(_03921_),
    .B2(_03923_),
    .ZN(_03924_));
 INV_X1 _27261_ (.A(_22016_),
    .ZN(_03925_));
 INV_X1 _27262_ (.A(_22017_),
    .ZN(_03926_));
 OAI21_X1 _27263_ (.A(_03925_),
    .B1(_03903_),
    .B2(_03926_),
    .ZN(_03927_));
 OAI21_X2 _27264_ (.A(_03919_),
    .B1(_03924_),
    .B2(_03927_),
    .ZN(_03928_));
 AOI21_X2 _27265_ (.A(_03918_),
    .B1(_03894_),
    .B2(_03928_),
    .ZN(_03929_));
 BUF_X4 _27266_ (.A(_03929_),
    .Z(_03930_));
 CLKBUF_X3 _27267_ (.A(_03930_),
    .Z(_03931_));
 MUX2_X2 _27268_ (.A(\g_reduce0[0].adder.x[10] ),
    .B(\g_reduce0[2].adder.x[10] ),
    .S(_03931_),
    .Z(_22119_));
 MUX2_X2 _27269_ (.A(_21997_),
    .B(_00565_),
    .S(_03931_),
    .Z(_14159_));
 BUF_X1 _27270_ (.A(_22032_),
    .Z(_03932_));
 NAND2_X1 _27271_ (.A1(_03887_),
    .A2(_03932_),
    .ZN(_03933_));
 MUX2_X2 _27272_ (.A(_00572_),
    .B(_22006_),
    .S(_03930_),
    .Z(_03934_));
 CLKBUF_X3 _27273_ (.A(_03931_),
    .Z(_03935_));
 MUX2_X1 _27274_ (.A(_00571_),
    .B(_22003_),
    .S(_03935_),
    .Z(_03936_));
 MUX2_X1 _27275_ (.A(_03934_),
    .B(_03936_),
    .S(_03887_),
    .Z(_03937_));
 INV_X1 _27276_ (.A(_03937_),
    .ZN(_03938_));
 BUF_X1 _27277_ (.A(_03932_),
    .Z(_03939_));
 OAI21_X2 _27278_ (.A(_03933_),
    .B1(_03938_),
    .B2(_03939_),
    .ZN(_03940_));
 CLKBUF_X2 _27279_ (.A(_22031_),
    .Z(_03941_));
 NOR2_X1 _27280_ (.A1(\g_reduce0[2].adder.x[11] ),
    .A2(_21997_),
    .ZN(_03942_));
 NOR2_X1 _27281_ (.A1(_03941_),
    .A2(_03942_),
    .ZN(_03943_));
 NOR2_X1 _27282_ (.A1(\g_reduce0[0].adder.x[11] ),
    .A2(_00565_),
    .ZN(_03944_));
 NOR2_X1 _27283_ (.A1(_03941_),
    .A2(_03944_),
    .ZN(_03945_));
 MUX2_X2 _27284_ (.A(_03943_),
    .B(_03945_),
    .S(_03929_),
    .Z(_03946_));
 XNOR2_X2 _27285_ (.A(_03881_),
    .B(_03946_),
    .ZN(_03947_));
 NOR2_X1 _27286_ (.A1(\g_reduce0[0].adder.x[13] ),
    .A2(_00573_),
    .ZN(_03948_));
 NOR2_X1 _27287_ (.A1(\g_reduce0[2].adder.x[13] ),
    .A2(_21991_),
    .ZN(_03949_));
 MUX2_X1 _27288_ (.A(_03948_),
    .B(_03949_),
    .S(_03908_),
    .Z(_03950_));
 NOR2_X2 _27289_ (.A1(\g_reduce0[0].adder.x[12] ),
    .A2(_00570_),
    .ZN(_03951_));
 INV_X1 _27290_ (.A(_03951_),
    .ZN(_03952_));
 NAND2_X1 _27291_ (.A1(_03916_),
    .A2(_03952_),
    .ZN(_03953_));
 AOI211_X2 _27292_ (.A(_03918_),
    .B(_03953_),
    .C1(_03928_),
    .C2(_03894_),
    .ZN(_03954_));
 NOR2_X2 _27293_ (.A1(\g_reduce0[2].adder.x[12] ),
    .A2(_21994_),
    .ZN(_03955_));
 NOR2_X1 _27294_ (.A1(_03881_),
    .A2(_03955_),
    .ZN(_03956_));
 AOI211_X2 _27295_ (.A(_03911_),
    .B(_03954_),
    .C1(_03956_),
    .C2(_03907_),
    .ZN(_03957_));
 OAI21_X1 _27296_ (.A(_03876_),
    .B1(_03950_),
    .B2(_03957_),
    .ZN(_03958_));
 OR3_X1 _27297_ (.A1(_03876_),
    .A2(_03950_),
    .A3(_03957_),
    .ZN(_03959_));
 MUX2_X2 _27298_ (.A(_03951_),
    .B(_03955_),
    .S(_03907_),
    .Z(_03960_));
 INV_X1 _27299_ (.A(\g_reduce0[2].adder.x[10] ),
    .ZN(_03961_));
 NAND2_X1 _27300_ (.A1(\g_reduce0[0].adder.x[10] ),
    .A2(_03961_),
    .ZN(_03962_));
 AOI211_X2 _27301_ (.A(_03918_),
    .B(_03962_),
    .C1(_03928_),
    .C2(_03894_),
    .ZN(_03963_));
 NOR2_X1 _27302_ (.A1(\g_reduce0[0].adder.x[10] ),
    .A2(_03961_),
    .ZN(_03964_));
 INV_X1 _27303_ (.A(_03964_),
    .ZN(_03965_));
 NOR3_X2 _27304_ (.A1(_03906_),
    .A2(_03895_),
    .A3(_03965_),
    .ZN(_03966_));
 INV_X1 _27305_ (.A(_03888_),
    .ZN(_03967_));
 OAI21_X2 _27306_ (.A(_03967_),
    .B1(_03885_),
    .B2(_03965_),
    .ZN(_03968_));
 NOR3_X4 _27307_ (.A1(_03963_),
    .A2(_03966_),
    .A3(_03968_),
    .ZN(_03969_));
 AND2_X1 _27308_ (.A1(_03881_),
    .A2(_03942_),
    .ZN(_03970_));
 AND2_X1 _27309_ (.A1(_03881_),
    .A2(_03944_),
    .ZN(_03971_));
 MUX2_X2 _27310_ (.A(_03970_),
    .B(_03971_),
    .S(_03930_),
    .Z(_03972_));
 NOR3_X4 _27311_ (.A1(_03960_),
    .A2(_03969_),
    .A3(_03972_),
    .ZN(_03973_));
 AOI221_X2 _27312_ (.A(_03947_),
    .B1(_03958_),
    .B2(_03959_),
    .C1(_03973_),
    .C2(_03911_),
    .ZN(_03974_));
 OAI21_X2 _27313_ (.A(_03974_),
    .B1(_03973_),
    .B2(_03911_),
    .ZN(_03975_));
 NOR2_X1 _27314_ (.A1(_03948_),
    .A2(_03951_),
    .ZN(_03976_));
 AND2_X1 _27315_ (.A1(_03930_),
    .A2(_03976_),
    .ZN(_03977_));
 NOR2_X1 _27316_ (.A1(_03949_),
    .A2(_03955_),
    .ZN(_03978_));
 AND2_X1 _27317_ (.A1(_03908_),
    .A2(_03978_),
    .ZN(_03979_));
 OAI221_X2 _27318_ (.A(_03910_),
    .B1(_03916_),
    .B2(_03946_),
    .C1(_03977_),
    .C2(_03979_),
    .ZN(_03980_));
 NAND2_X1 _27319_ (.A1(_03876_),
    .A2(_03950_),
    .ZN(_03981_));
 AOI211_X2 _27320_ (.A(_03911_),
    .B(_03973_),
    .C1(_03980_),
    .C2(_03981_),
    .ZN(_03982_));
 AOI211_X2 _27321_ (.A(_03960_),
    .B(_03972_),
    .C1(_03969_),
    .C2(_03941_),
    .ZN(_03983_));
 NAND2_X1 _27322_ (.A1(_03876_),
    .A2(_03911_),
    .ZN(_03984_));
 NAND2_X1 _27323_ (.A1(_03910_),
    .A2(_03911_),
    .ZN(_03985_));
 INV_X1 _27324_ (.A(_03948_),
    .ZN(_03986_));
 INV_X1 _27325_ (.A(_03949_),
    .ZN(_03987_));
 MUX2_X2 _27326_ (.A(_03986_),
    .B(_03987_),
    .S(_03907_),
    .Z(_03988_));
 MUX2_X1 _27327_ (.A(_03984_),
    .B(_03985_),
    .S(_03988_),
    .Z(_03989_));
 INV_X1 _27328_ (.A(_03955_),
    .ZN(_03990_));
 MUX2_X2 _27329_ (.A(_03952_),
    .B(_03990_),
    .S(_03908_),
    .Z(_03991_));
 OR3_X2 _27330_ (.A1(_03963_),
    .A2(_03966_),
    .A3(_03968_),
    .ZN(_03992_));
 NAND2_X1 _27331_ (.A1(_03881_),
    .A2(_03942_),
    .ZN(_03993_));
 NAND2_X1 _27332_ (.A1(_03881_),
    .A2(_03944_),
    .ZN(_03994_));
 MUX2_X2 _27333_ (.A(_03993_),
    .B(_03994_),
    .S(_03930_),
    .Z(_03995_));
 NAND3_X4 _27334_ (.A1(_03991_),
    .A2(_03992_),
    .A3(_03995_),
    .ZN(_03996_));
 OAI22_X4 _27335_ (.A1(_03884_),
    .A2(_03983_),
    .B1(_03989_),
    .B2(_03996_),
    .ZN(_03997_));
 NOR2_X4 _27336_ (.A1(_03982_),
    .A2(_03997_),
    .ZN(_03998_));
 MUX2_X1 _27337_ (.A(_00564_),
    .B(_22024_),
    .S(_03931_),
    .Z(_03999_));
 MUX2_X1 _27338_ (.A(_00563_),
    .B(_22021_),
    .S(_03935_),
    .Z(_04000_));
 MUX2_X1 _27339_ (.A(_03999_),
    .B(_04000_),
    .S(_03887_),
    .Z(_04001_));
 MUX2_X1 _27340_ (.A(_00561_),
    .B(_00562_),
    .S(_03935_),
    .Z(_04002_));
 MUX2_X1 _27341_ (.A(_00560_),
    .B(_22027_),
    .S(_03935_),
    .Z(_04003_));
 MUX2_X1 _27342_ (.A(_04002_),
    .B(_04003_),
    .S(_03887_),
    .Z(_04004_));
 INV_X1 _27343_ (.A(_03939_),
    .ZN(_04005_));
 MUX2_X1 _27344_ (.A(_04001_),
    .B(_04004_),
    .S(_04005_),
    .Z(_04006_));
 MUX2_X1 _27345_ (.A(_00569_),
    .B(_22012_),
    .S(_03935_),
    .Z(_04007_));
 MUX2_X1 _27346_ (.A(_00568_),
    .B(_22009_),
    .S(_03935_),
    .Z(_04008_));
 MUX2_X1 _27347_ (.A(_04007_),
    .B(_04008_),
    .S(_03887_),
    .Z(_04009_));
 MUX2_X1 _27348_ (.A(_00567_),
    .B(_22018_),
    .S(_03935_),
    .Z(_04010_));
 MUX2_X1 _27349_ (.A(_00566_),
    .B(_22015_),
    .S(_03935_),
    .Z(_04011_));
 MUX2_X1 _27350_ (.A(_04010_),
    .B(_04011_),
    .S(_03887_),
    .Z(_04012_));
 MUX2_X1 _27351_ (.A(_04009_),
    .B(_04012_),
    .S(_04005_),
    .Z(_04013_));
 MUX2_X1 _27352_ (.A(_04006_),
    .B(_04013_),
    .S(_03947_),
    .Z(_04014_));
 OAI22_X2 _27353_ (.A1(_03940_),
    .A2(_03975_),
    .B1(_03998_),
    .B2(_04014_),
    .ZN(_22096_));
 MUX2_X1 _27354_ (.A(_03999_),
    .B(_04010_),
    .S(_03939_),
    .Z(_04015_));
 MUX2_X1 _27355_ (.A(_04000_),
    .B(_04003_),
    .S(_04005_),
    .Z(_04016_));
 CLKBUF_X3 _27356_ (.A(_03886_),
    .Z(_04017_));
 MUX2_X1 _27357_ (.A(_04015_),
    .B(_04016_),
    .S(_04017_),
    .Z(_04018_));
 MUX2_X1 _27358_ (.A(_04008_),
    .B(_04011_),
    .S(_04005_),
    .Z(_04019_));
 MUX2_X1 _27359_ (.A(_03934_),
    .B(_04007_),
    .S(_04005_),
    .Z(_04020_));
 MUX2_X1 _27360_ (.A(_04019_),
    .B(_04020_),
    .S(_03887_),
    .Z(_04021_));
 MUX2_X1 _27361_ (.A(_04018_),
    .B(_04021_),
    .S(_03947_),
    .Z(_04022_));
 NOR2_X1 _27362_ (.A1(_03998_),
    .A2(_04022_),
    .ZN(_04023_));
 AOI21_X2 _27363_ (.A(_03939_),
    .B1(_03936_),
    .B2(_04017_),
    .ZN(_04024_));
 INV_X1 _27364_ (.A(_03975_),
    .ZN(_04025_));
 AOI21_X2 _27365_ (.A(_04023_),
    .B1(_04024_),
    .B2(_04025_),
    .ZN(_14153_));
 INV_X1 _27366_ (.A(_14153_),
    .ZN(_14149_));
 INV_X1 _27367_ (.A(_22096_),
    .ZN(_22099_));
 NOR2_X1 _27368_ (.A1(_03947_),
    .A2(_03998_),
    .ZN(_04026_));
 NAND2_X1 _27369_ (.A1(_04024_),
    .A2(_04026_),
    .ZN(_22052_));
 INV_X1 _27370_ (.A(_22052_),
    .ZN(_22055_));
 OR3_X1 _27371_ (.A1(_03940_),
    .A2(_03947_),
    .A3(_03998_),
    .ZN(_22045_));
 INV_X1 _27372_ (.A(_22045_),
    .ZN(_22048_));
 MUX2_X1 _27373_ (.A(_00568_),
    .B(_00571_),
    .S(_03939_),
    .Z(_04027_));
 MUX2_X1 _27374_ (.A(_22009_),
    .B(_22003_),
    .S(_03939_),
    .Z(_04028_));
 MUX2_X1 _27375_ (.A(_04027_),
    .B(_04028_),
    .S(_03931_),
    .Z(_04029_));
 NOR2_X1 _27376_ (.A1(_04017_),
    .A2(_03939_),
    .ZN(_04030_));
 AOI22_X2 _27377_ (.A1(_04017_),
    .A2(_04029_),
    .B1(_04030_),
    .B2(_03934_),
    .ZN(_04031_));
 NAND2_X1 _27378_ (.A1(_04026_),
    .A2(_04031_),
    .ZN(_22079_));
 INV_X1 _27379_ (.A(_22079_),
    .ZN(_22083_));
 MUX2_X1 _27380_ (.A(_03937_),
    .B(_04009_),
    .S(_04005_),
    .Z(_04032_));
 NAND2_X1 _27381_ (.A1(_04017_),
    .A2(_04005_),
    .ZN(_04033_));
 MUX2_X1 _27382_ (.A(_04032_),
    .B(_04033_),
    .S(_03947_),
    .Z(_04034_));
 OR2_X1 _27383_ (.A1(_03998_),
    .A2(_04034_),
    .ZN(_22059_));
 INV_X1 _27384_ (.A(_22059_),
    .ZN(_22062_));
 INV_X1 _27385_ (.A(_04024_),
    .ZN(_04035_));
 XNOR2_X2 _27386_ (.A(_03916_),
    .B(_03946_),
    .ZN(_04036_));
 MUX2_X1 _27387_ (.A(_04035_),
    .B(_04021_),
    .S(_04036_),
    .Z(_04037_));
 NOR2_X1 _27388_ (.A1(_03998_),
    .A2(_04037_),
    .ZN(_22066_));
 INV_X1 _27389_ (.A(_22066_),
    .ZN(_22069_));
 MUX2_X1 _27390_ (.A(_03940_),
    .B(_04013_),
    .S(_04036_),
    .Z(_04038_));
 NOR2_X1 _27391_ (.A1(_03998_),
    .A2(_04038_),
    .ZN(_22073_));
 INV_X1 _27392_ (.A(_22073_),
    .ZN(_22076_));
 MUX2_X1 _27393_ (.A(_22018_),
    .B(_22012_),
    .S(_03932_),
    .Z(_04039_));
 MUX2_X1 _27394_ (.A(_22021_),
    .B(_22015_),
    .S(_03932_),
    .Z(_04040_));
 MUX2_X1 _27395_ (.A(_04039_),
    .B(_04040_),
    .S(_03886_),
    .Z(_04041_));
 MUX2_X1 _27396_ (.A(_00567_),
    .B(_00569_),
    .S(_03932_),
    .Z(_04042_));
 MUX2_X1 _27397_ (.A(_00563_),
    .B(_00566_),
    .S(_03932_),
    .Z(_04043_));
 MUX2_X1 _27398_ (.A(_04042_),
    .B(_04043_),
    .S(_03886_),
    .Z(_04044_));
 MUX2_X1 _27399_ (.A(_04041_),
    .B(_04044_),
    .S(_03908_),
    .Z(_04045_));
 NOR2_X1 _27400_ (.A1(_03947_),
    .A2(_04045_),
    .ZN(_04046_));
 AOI21_X1 _27401_ (.A(_04046_),
    .B1(_04031_),
    .B2(_03947_),
    .ZN(_04047_));
 NOR2_X1 _27402_ (.A1(_03998_),
    .A2(_04047_),
    .ZN(_22090_));
 INV_X1 _27403_ (.A(_22090_),
    .ZN(_22093_));
 MUX2_X1 _27404_ (.A(_04001_),
    .B(_04012_),
    .S(_03939_),
    .Z(_04048_));
 MUX2_X1 _27405_ (.A(_04032_),
    .B(_04048_),
    .S(_04036_),
    .Z(_04049_));
 OAI22_X2 _27406_ (.A1(_03975_),
    .A2(_04033_),
    .B1(_04049_),
    .B2(_03998_),
    .ZN(_22040_));
 INV_X1 _27407_ (.A(_22040_),
    .ZN(_22086_));
 XOR2_X2 _27408_ (.A(\g_reduce0[0].adder.x[15] ),
    .B(\g_reduce0[2].adder.x[15] ),
    .Z(_04050_));
 CLKBUF_X3 _27409_ (.A(_04050_),
    .Z(_04051_));
 BUF_X2 _27410_ (.A(_22054_),
    .Z(_04052_));
 BUF_X2 _27411_ (.A(_22047_),
    .Z(_04053_));
 INV_X1 _27412_ (.A(_04053_),
    .ZN(_04054_));
 BUF_X2 _27413_ (.A(_22082_),
    .Z(_04055_));
 CLKBUF_X3 _27414_ (.A(_22061_),
    .Z(_04056_));
 INV_X1 _27415_ (.A(_22067_),
    .ZN(_04057_));
 BUF_X4 _27416_ (.A(_22075_),
    .Z(_04058_));
 OAI21_X1 _27417_ (.A(_22068_),
    .B1(_04058_),
    .B2(_22074_),
    .ZN(_04059_));
 AOI21_X1 _27418_ (.A(_04056_),
    .B1(_04057_),
    .B2(_04059_),
    .ZN(_04060_));
 NOR2_X1 _27419_ (.A1(_22063_),
    .A2(_04060_),
    .ZN(_04061_));
 INV_X1 _27420_ (.A(_22063_),
    .ZN(_04062_));
 NOR2_X1 _27421_ (.A1(_22074_),
    .A2(_22091_),
    .ZN(_04063_));
 NAND3_X1 _27422_ (.A1(_04062_),
    .A2(_04057_),
    .A3(_04063_),
    .ZN(_04064_));
 INV_X1 _27423_ (.A(_22042_),
    .ZN(_04065_));
 INV_X1 _27424_ (.A(_22043_),
    .ZN(_04066_));
 AOI21_X1 _27425_ (.A(_22036_),
    .B1(_14150_),
    .B2(_22037_),
    .ZN(_04067_));
 OAI21_X1 _27426_ (.A(_04065_),
    .B1(_04066_),
    .B2(_04067_),
    .ZN(_04068_));
 BUF_X2 _27427_ (.A(_22092_),
    .Z(_04069_));
 AOI21_X1 _27428_ (.A(_04064_),
    .B1(_04068_),
    .B2(_04069_),
    .ZN(_04070_));
 NOR3_X1 _27429_ (.A1(_04055_),
    .A2(_04061_),
    .A3(_04070_),
    .ZN(_04071_));
 OAI21_X1 _27430_ (.A(_04054_),
    .B1(_04071_),
    .B2(_22084_),
    .ZN(_04072_));
 INV_X1 _27431_ (.A(_22049_),
    .ZN(_04073_));
 AOI21_X1 _27432_ (.A(_04052_),
    .B1(_04072_),
    .B2(_04073_),
    .ZN(_04074_));
 NOR2_X1 _27433_ (.A1(_22056_),
    .A2(_04074_),
    .ZN(_04075_));
 NOR2_X1 _27434_ (.A1(_04051_),
    .A2(_04075_),
    .ZN(_04076_));
 XNOR2_X1 _27435_ (.A(\g_reduce0[0].adder.x[15] ),
    .B(\g_reduce0[2].adder.x[15] ),
    .ZN(_04077_));
 CLKBUF_X3 _27436_ (.A(_04077_),
    .Z(_04078_));
 CLKBUF_X3 _27437_ (.A(_04078_),
    .Z(_04079_));
 NOR2_X1 _27438_ (.A1(_04053_),
    .A2(_22046_),
    .ZN(_04080_));
 NOR2_X1 _27439_ (.A1(_22081_),
    .A2(_22046_),
    .ZN(_04081_));
 INV_X1 _27440_ (.A(_04055_),
    .ZN(_04082_));
 INV_X1 _27441_ (.A(_22077_),
    .ZN(_04083_));
 AOI21_X4 _27442_ (.A(_22068_),
    .B1(_04058_),
    .B2(_04083_),
    .ZN(_04084_));
 OR2_X1 _27443_ (.A1(_22070_),
    .A2(_22060_),
    .ZN(_04085_));
 OAI22_X4 _27444_ (.A1(_04056_),
    .A2(_22060_),
    .B1(_04084_),
    .B2(_04085_),
    .ZN(_04086_));
 OR3_X1 _27445_ (.A1(_22077_),
    .A2(_22094_),
    .A3(_04085_),
    .ZN(_04087_));
 INV_X1 _27446_ (.A(_22087_),
    .ZN(_04088_));
 INV_X1 _27447_ (.A(_22088_),
    .ZN(_04089_));
 AOI21_X1 _27448_ (.A(_22038_),
    .B1(_14154_),
    .B2(_22039_),
    .ZN(_04090_));
 OAI21_X2 _27449_ (.A(_04088_),
    .B1(_04089_),
    .B2(_04090_),
    .ZN(_04091_));
 INV_X1 _27450_ (.A(_04069_),
    .ZN(_04092_));
 AOI21_X2 _27451_ (.A(_04087_),
    .B1(_04091_),
    .B2(_04092_),
    .ZN(_04093_));
 OR3_X1 _27452_ (.A1(_04082_),
    .A2(_04086_),
    .A3(_04093_),
    .ZN(_04094_));
 AOI21_X1 _27453_ (.A(_04080_),
    .B1(_04081_),
    .B2(_04094_),
    .ZN(_04095_));
 AOI21_X1 _27454_ (.A(_22053_),
    .B1(_04095_),
    .B2(_04052_),
    .ZN(_04096_));
 OR2_X1 _27455_ (.A1(_04079_),
    .A2(_04096_),
    .ZN(_04097_));
 NAND4_X1 _27456_ (.A1(_04017_),
    .A2(_04005_),
    .A3(_04036_),
    .A4(_04097_),
    .ZN(_04098_));
 INV_X1 _27457_ (.A(_03941_),
    .ZN(_04099_));
 OAI211_X2 _27458_ (.A(_03991_),
    .B(_03995_),
    .C1(_03992_),
    .C2(_04099_),
    .ZN(_04100_));
 NOR2_X1 _27459_ (.A1(_03910_),
    .A2(_03883_),
    .ZN(_04101_));
 NOR2_X1 _27460_ (.A1(_03876_),
    .A2(_03883_),
    .ZN(_04102_));
 MUX2_X1 _27461_ (.A(_04101_),
    .B(_04102_),
    .S(_03988_),
    .Z(_04103_));
 AOI22_X4 _27462_ (.A1(_03912_),
    .A2(_04100_),
    .B1(_04103_),
    .B2(_03973_),
    .ZN(_04104_));
 OR2_X1 _27463_ (.A1(_03941_),
    .A2(_03942_),
    .ZN(_04105_));
 OR2_X1 _27464_ (.A1(_03941_),
    .A2(_03944_),
    .ZN(_04106_));
 MUX2_X1 _27465_ (.A(_04105_),
    .B(_04106_),
    .S(_03930_),
    .Z(_04107_));
 NAND2_X1 _27466_ (.A1(_03930_),
    .A2(_03976_),
    .ZN(_04108_));
 NAND2_X1 _27467_ (.A1(_03908_),
    .A2(_03978_),
    .ZN(_04109_));
 AOI221_X2 _27468_ (.A(_03876_),
    .B1(_03881_),
    .B2(_04107_),
    .C1(_04108_),
    .C2(_04109_),
    .ZN(_04110_));
 NOR2_X1 _27469_ (.A1(_03910_),
    .A2(_03988_),
    .ZN(_04111_));
 OAI211_X4 _27470_ (.A(_03883_),
    .B(_03996_),
    .C1(_04110_),
    .C2(_04111_),
    .ZN(_04112_));
 AOI21_X2 _27471_ (.A(_04098_),
    .B1(_04104_),
    .B2(_04112_),
    .ZN(_04113_));
 NOR2_X1 _27472_ (.A1(_04076_),
    .A2(_04113_),
    .ZN(_04114_));
 BUF_X4 _27473_ (.A(_04114_),
    .Z(_04115_));
 OR2_X1 _27474_ (.A1(_03947_),
    .A2(_04033_),
    .ZN(_04116_));
 AOI21_X4 _27475_ (.A(_04116_),
    .B1(_04104_),
    .B2(_04112_),
    .ZN(_04117_));
 AOI21_X1 _27476_ (.A(_04052_),
    .B1(_22053_),
    .B2(_04051_),
    .ZN(_04118_));
 NAND2_X1 _27477_ (.A1(_04073_),
    .A2(_04079_),
    .ZN(_04119_));
 OR2_X1 _27478_ (.A1(_04056_),
    .A2(_04055_),
    .ZN(_04120_));
 OAI22_X2 _27479_ (.A1(_04062_),
    .A2(_04055_),
    .B1(_04057_),
    .B2(_04120_),
    .ZN(_04121_));
 NOR2_X1 _27480_ (.A1(_04059_),
    .A2(_04120_),
    .ZN(_04122_));
 AOI21_X1 _27481_ (.A(_22042_),
    .B1(_14151_),
    .B2(_22043_),
    .ZN(_04123_));
 OAI21_X1 _27482_ (.A(_04063_),
    .B1(_04123_),
    .B2(_04092_),
    .ZN(_04124_));
 AOI211_X2 _27483_ (.A(_22084_),
    .B(_04121_),
    .C1(_04122_),
    .C2(_04124_),
    .ZN(_04125_));
 NOR2_X1 _27484_ (.A1(_04053_),
    .A2(_04125_),
    .ZN(_04126_));
 OAI21_X1 _27485_ (.A(_04118_),
    .B1(_04119_),
    .B2(_04126_),
    .ZN(_04127_));
 AOI21_X1 _27486_ (.A(_22081_),
    .B1(_22060_),
    .B2(_04055_),
    .ZN(_04128_));
 NAND2_X1 _27487_ (.A1(_04056_),
    .A2(_04055_),
    .ZN(_04129_));
 NOR2_X1 _27488_ (.A1(_22077_),
    .A2(_22094_),
    .ZN(_04130_));
 AOI21_X1 _27489_ (.A(_22087_),
    .B1(_14155_),
    .B2(_22088_),
    .ZN(_04131_));
 OAI21_X1 _27490_ (.A(_04130_),
    .B1(_04131_),
    .B2(_04069_),
    .ZN(_04132_));
 AOI21_X2 _27491_ (.A(_22070_),
    .B1(_04084_),
    .B2(_04132_),
    .ZN(_04133_));
 OAI21_X1 _27492_ (.A(_04128_),
    .B1(_04129_),
    .B2(_04133_),
    .ZN(_04134_));
 NAND2_X1 _27493_ (.A1(_04053_),
    .A2(_04134_),
    .ZN(_04135_));
 NOR3_X1 _27494_ (.A1(_22053_),
    .A2(_22046_),
    .A3(_04079_),
    .ZN(_04136_));
 AOI22_X2 _27495_ (.A1(_22056_),
    .A2(_04079_),
    .B1(_04135_),
    .B2(_04136_),
    .ZN(_04137_));
 AND2_X2 _27496_ (.A1(_04127_),
    .A2(_04137_),
    .ZN(_04138_));
 XNOR2_X2 _27497_ (.A(_04117_),
    .B(_04138_),
    .ZN(_04139_));
 BUF_X2 _27498_ (.A(_04139_),
    .Z(_04140_));
 NAND2_X1 _27499_ (.A1(_04054_),
    .A2(_04077_),
    .ZN(_04141_));
 OR4_X1 _27500_ (.A1(_04055_),
    .A2(_04061_),
    .A3(_04070_),
    .A4(_04141_),
    .ZN(_04142_));
 AND2_X1 _27501_ (.A1(_04050_),
    .A2(_04081_),
    .ZN(_04143_));
 OAI21_X2 _27502_ (.A(_04143_),
    .B1(_04093_),
    .B2(_04086_),
    .ZN(_04144_));
 AOI22_X2 _27503_ (.A1(_04050_),
    .A2(_04080_),
    .B1(_04143_),
    .B2(_04082_),
    .ZN(_04145_));
 AOI21_X1 _27504_ (.A(_22049_),
    .B1(_04054_),
    .B2(_22084_),
    .ZN(_04146_));
 OR2_X1 _27505_ (.A1(_04050_),
    .A2(_04146_),
    .ZN(_04147_));
 NAND4_X4 _27506_ (.A1(_04142_),
    .A2(_04144_),
    .A3(_04145_),
    .A4(_04147_),
    .ZN(_04148_));
 XOR2_X2 _27507_ (.A(_04052_),
    .B(_04148_),
    .Z(_04149_));
 OR2_X1 _27508_ (.A1(_04050_),
    .A2(_04125_),
    .ZN(_04150_));
 OAI21_X2 _27509_ (.A(_04150_),
    .B1(_04134_),
    .B2(_04078_),
    .ZN(_04151_));
 XNOR2_X2 _27510_ (.A(_04053_),
    .B(_04151_),
    .ZN(_04152_));
 NOR3_X1 _27511_ (.A1(_04079_),
    .A2(_04086_),
    .A3(_04093_),
    .ZN(_04153_));
 OR2_X1 _27512_ (.A1(_04061_),
    .A2(_04070_),
    .ZN(_04154_));
 AOI21_X2 _27513_ (.A(_04153_),
    .B1(_04154_),
    .B2(_04079_),
    .ZN(_04155_));
 XNOR2_X2 _27514_ (.A(_04055_),
    .B(_04155_),
    .ZN(_04156_));
 INV_X1 _27515_ (.A(_04059_),
    .ZN(_04157_));
 AOI21_X1 _27516_ (.A(_22067_),
    .B1(_04157_),
    .B2(_04124_),
    .ZN(_04158_));
 NOR2_X1 _27517_ (.A1(_04050_),
    .A2(_04158_),
    .ZN(_04159_));
 AOI21_X4 _27518_ (.A(_04159_),
    .B1(_04133_),
    .B2(_04050_),
    .ZN(_04160_));
 XNOR2_X2 _27519_ (.A(_04056_),
    .B(_04160_),
    .ZN(_04161_));
 INV_X1 _27520_ (.A(_22068_),
    .ZN(_04162_));
 AND2_X1 _27521_ (.A1(_04069_),
    .A2(_04068_),
    .ZN(_04163_));
 OR2_X1 _27522_ (.A1(_22074_),
    .A2(_22091_),
    .ZN(_04164_));
 OAI221_X2 _27523_ (.A(_04078_),
    .B1(_04163_),
    .B2(_04164_),
    .C1(_22074_),
    .C2(_04058_),
    .ZN(_04165_));
 NOR2_X1 _27524_ (.A1(_22077_),
    .A2(_04078_),
    .ZN(_04166_));
 AOI21_X1 _27525_ (.A(_22094_),
    .B1(_04091_),
    .B2(_04092_),
    .ZN(_04167_));
 OAI21_X2 _27526_ (.A(_04166_),
    .B1(_04167_),
    .B2(_04058_),
    .ZN(_04168_));
 AND3_X1 _27527_ (.A1(_04162_),
    .A2(_04165_),
    .A3(_04168_),
    .ZN(_04169_));
 AOI21_X4 _27528_ (.A(_04162_),
    .B1(_04165_),
    .B2(_04168_),
    .ZN(_04170_));
 NOR2_X1 _27529_ (.A1(_04092_),
    .A2(_04123_),
    .ZN(_04171_));
 OAI21_X1 _27530_ (.A(_04078_),
    .B1(_04171_),
    .B2(_22091_),
    .ZN(_04172_));
 INV_X1 _27531_ (.A(_22094_),
    .ZN(_04173_));
 OAI21_X1 _27532_ (.A(_04173_),
    .B1(_04131_),
    .B2(_04069_),
    .ZN(_04174_));
 OAI21_X2 _27533_ (.A(_04172_),
    .B1(_04174_),
    .B2(_04078_),
    .ZN(_04175_));
 XOR2_X2 _27534_ (.A(_04058_),
    .B(_04175_),
    .Z(_04176_));
 XOR2_X1 _27535_ (.A(_14151_),
    .B(_22043_),
    .Z(_04177_));
 NAND2_X1 _27536_ (.A1(_04078_),
    .A2(_04177_),
    .ZN(_04178_));
 XOR2_X1 _27537_ (.A(_14155_),
    .B(_22088_),
    .Z(_04179_));
 NAND2_X1 _27538_ (.A1(_04051_),
    .A2(_04179_),
    .ZN(_04180_));
 NAND2_X1 _27539_ (.A1(_04178_),
    .A2(_04180_),
    .ZN(_04181_));
 MUX2_X2 _27540_ (.A(_14156_),
    .B(_14152_),
    .S(_04079_),
    .Z(_04182_));
 NOR2_X1 _27541_ (.A1(_04181_),
    .A2(_04182_),
    .ZN(_04183_));
 AND2_X1 _27542_ (.A1(_04078_),
    .A2(_04068_),
    .ZN(_04184_));
 NOR2_X1 _27543_ (.A1(_04078_),
    .A2(_04091_),
    .ZN(_04185_));
 OAI21_X2 _27544_ (.A(_04069_),
    .B1(_04184_),
    .B2(_04185_),
    .ZN(_04186_));
 OR3_X2 _27545_ (.A1(_04069_),
    .A2(_04184_),
    .A3(_04185_),
    .ZN(_04187_));
 AOI21_X2 _27546_ (.A(_04183_),
    .B1(_04186_),
    .B2(_04187_),
    .ZN(_04188_));
 OAI22_X4 _27547_ (.A1(_04169_),
    .A2(_04170_),
    .B1(_04176_),
    .B2(_04188_),
    .ZN(_04189_));
 AOI21_X4 _27548_ (.A(_04156_),
    .B1(_04161_),
    .B2(_04189_),
    .ZN(_04190_));
 OAI21_X4 _27549_ (.A(_04149_),
    .B1(_04152_),
    .B2(_04190_),
    .ZN(_04191_));
 AND2_X1 _27550_ (.A1(_03931_),
    .A2(_04041_),
    .ZN(_04192_));
 AOI21_X1 _27551_ (.A(_04192_),
    .B1(_04044_),
    .B2(_03908_),
    .ZN(_04193_));
 OR3_X1 _27552_ (.A1(_00561_),
    .A2(_03886_),
    .A3(_03939_),
    .ZN(_04194_));
 OR3_X1 _27553_ (.A1(_00562_),
    .A2(_04017_),
    .A3(_03939_),
    .ZN(_04195_));
 MUX2_X1 _27554_ (.A(_04194_),
    .B(_04195_),
    .S(_03931_),
    .Z(_04196_));
 INV_X1 _27555_ (.A(_00560_),
    .ZN(_04197_));
 NAND2_X1 _27556_ (.A1(_04197_),
    .A2(_04017_),
    .ZN(_04198_));
 INV_X1 _27557_ (.A(_22027_),
    .ZN(_04199_));
 NAND2_X1 _27558_ (.A1(_04199_),
    .A2(_04017_),
    .ZN(_04200_));
 MUX2_X1 _27559_ (.A(_04198_),
    .B(_04200_),
    .S(_03931_),
    .Z(_04201_));
 OAI221_X1 _27560_ (.A(_04196_),
    .B1(_04201_),
    .B2(_04005_),
    .C1(_03933_),
    .C2(_03999_),
    .ZN(_04202_));
 MUX2_X1 _27561_ (.A(_04193_),
    .B(_04202_),
    .S(_04036_),
    .Z(_04203_));
 XOR2_X2 _27562_ (.A(_04056_),
    .B(_04160_),
    .Z(_04204_));
 AND2_X1 _27563_ (.A1(_04178_),
    .A2(_04180_),
    .ZN(_04205_));
 AND2_X1 _27564_ (.A1(_22098_),
    .A2(_04078_),
    .ZN(_04206_));
 AOI21_X4 _27565_ (.A(_04206_),
    .B1(_04051_),
    .B2(_22100_),
    .ZN(_04207_));
 NAND2_X1 _27566_ (.A1(_04205_),
    .A2(_04207_),
    .ZN(_04208_));
 NOR4_X4 _27567_ (.A1(_04152_),
    .A2(_04204_),
    .A3(_04176_),
    .A4(_04208_),
    .ZN(_04209_));
 AND2_X1 _27568_ (.A1(_04079_),
    .A2(_04209_),
    .ZN(_04210_));
 OAI211_X2 _27569_ (.A(_04203_),
    .B(_04210_),
    .C1(_03982_),
    .C2(_03997_),
    .ZN(_04211_));
 NAND2_X1 _27570_ (.A1(_04079_),
    .A2(_04209_),
    .ZN(_04212_));
 AOI222_X2 _27571_ (.A1(_03883_),
    .A2(_03996_),
    .B1(_04030_),
    .B2(_03934_),
    .C1(_04029_),
    .C2(_04017_),
    .ZN(_04213_));
 NAND2_X1 _27572_ (.A1(_03974_),
    .A2(_04213_),
    .ZN(_04214_));
 NOR3_X1 _27573_ (.A1(_00561_),
    .A2(_03886_),
    .A3(_03932_),
    .ZN(_04215_));
 NOR3_X1 _27574_ (.A1(_00562_),
    .A2(_03886_),
    .A3(_03932_),
    .ZN(_04216_));
 MUX2_X1 _27575_ (.A(_04215_),
    .B(_04216_),
    .S(_03930_),
    .Z(_04217_));
 NOR2_X1 _27576_ (.A1(_00560_),
    .A2(_03887_),
    .ZN(_04218_));
 NOR2_X1 _27577_ (.A1(_22027_),
    .A2(_03887_),
    .ZN(_04219_));
 MUX2_X1 _27578_ (.A(_04218_),
    .B(_04219_),
    .S(_03930_),
    .Z(_04220_));
 INV_X1 _27579_ (.A(_03933_),
    .ZN(_04221_));
 INV_X1 _27580_ (.A(_00564_),
    .ZN(_04222_));
 INV_X1 _27581_ (.A(_22024_),
    .ZN(_04223_));
 MUX2_X1 _27582_ (.A(_04222_),
    .B(_04223_),
    .S(_03930_),
    .Z(_04224_));
 AOI221_X2 _27583_ (.A(_04217_),
    .B1(_04220_),
    .B2(_03932_),
    .C1(_04221_),
    .C2(_04224_),
    .ZN(_04225_));
 MUX2_X1 _27584_ (.A(_04045_),
    .B(_04225_),
    .S(_04036_),
    .Z(_04226_));
 AOI21_X1 _27585_ (.A(_04226_),
    .B1(_04104_),
    .B2(_04112_),
    .ZN(_04227_));
 AND2_X1 _27586_ (.A1(_04051_),
    .A2(_04209_),
    .ZN(_04228_));
 OAI21_X1 _27587_ (.A(_04031_),
    .B1(_03973_),
    .B2(_03911_),
    .ZN(_04229_));
 NOR2_X1 _27588_ (.A1(_03881_),
    .A2(_03951_),
    .ZN(_04230_));
 MUX2_X1 _27589_ (.A(_03956_),
    .B(_04230_),
    .S(_03931_),
    .Z(_04231_));
 OAI22_X2 _27590_ (.A1(_03910_),
    .A2(_03988_),
    .B1(_04231_),
    .B2(_03884_),
    .ZN(_04232_));
 NOR3_X1 _27591_ (.A1(_03876_),
    .A2(_03950_),
    .A3(_03957_),
    .ZN(_04233_));
 OAI221_X2 _27592_ (.A(_04036_),
    .B1(_04232_),
    .B2(_04233_),
    .C1(_03996_),
    .C2(_03883_),
    .ZN(_04234_));
 OAI21_X1 _27593_ (.A(_04228_),
    .B1(_04229_),
    .B2(_04234_),
    .ZN(_04235_));
 OAI221_X1 _27594_ (.A(_04211_),
    .B1(_04212_),
    .B2(_04214_),
    .C1(_04227_),
    .C2(_04235_),
    .ZN(_04236_));
 OAI21_X1 _27595_ (.A(_04140_),
    .B1(_04191_),
    .B2(_04236_),
    .ZN(_04237_));
 NAND2_X2 _27596_ (.A1(_04115_),
    .A2(_04237_),
    .ZN(_22101_));
 INV_X1 _27597_ (.A(_22101_),
    .ZN(_22104_));
 XNOR2_X2 _27598_ (.A(_04054_),
    .B(_04151_),
    .ZN(_04238_));
 NAND2_X1 _27599_ (.A1(_04149_),
    .A2(_04238_),
    .ZN(_04239_));
 OR2_X1 _27600_ (.A1(_04169_),
    .A2(_04170_),
    .ZN(_04240_));
 XNOR2_X2 _27601_ (.A(_04058_),
    .B(_04175_),
    .ZN(_04241_));
 AND2_X1 _27602_ (.A1(_04187_),
    .A2(_04186_),
    .ZN(_04242_));
 NOR2_X2 _27603_ (.A1(_04242_),
    .A2(_04181_),
    .ZN(_04243_));
 AND3_X1 _27604_ (.A1(_04240_),
    .A2(_04241_),
    .A3(_04243_),
    .ZN(_04244_));
 NOR4_X2 _27605_ (.A1(_04156_),
    .A2(_04204_),
    .A3(_04239_),
    .A4(_04244_),
    .ZN(_04245_));
 NAND2_X2 _27606_ (.A1(_04127_),
    .A2(_04137_),
    .ZN(_04246_));
 OAI21_X1 _27607_ (.A(_04246_),
    .B1(_04075_),
    .B2(_04051_),
    .ZN(_04247_));
 OR2_X1 _27608_ (.A1(_04245_),
    .A2(_04247_),
    .ZN(_04248_));
 OR2_X1 _27609_ (.A1(_04097_),
    .A2(_04246_),
    .ZN(_04249_));
 OR2_X1 _27610_ (.A1(_04245_),
    .A2(_04249_),
    .ZN(_04250_));
 MUX2_X1 _27611_ (.A(_04248_),
    .B(_04250_),
    .S(_04117_),
    .Z(_04251_));
 XOR2_X2 _27612_ (.A(_22107_),
    .B(_04251_),
    .Z(_04252_));
 INV_X2 _27613_ (.A(_04252_),
    .ZN(_04253_));
 CLKBUF_X3 _27614_ (.A(_04253_),
    .Z(_22127_));
 INV_X1 _27615_ (.A(_04249_),
    .ZN(_04254_));
 INV_X1 _27616_ (.A(_04247_),
    .ZN(_04255_));
 NOR2_X1 _27617_ (.A1(_03947_),
    .A2(_04033_),
    .ZN(_04256_));
 OAI21_X2 _27618_ (.A(_04256_),
    .B1(_03997_),
    .B2(_03982_),
    .ZN(_04257_));
 MUX2_X1 _27619_ (.A(_04254_),
    .B(_04255_),
    .S(_04257_),
    .Z(_04258_));
 BUF_X4 _27620_ (.A(_04258_),
    .Z(_04259_));
 CLKBUF_X2 _27621_ (.A(_22103_),
    .Z(_04260_));
 INV_X2 _27622_ (.A(_04260_),
    .ZN(_04261_));
 MUX2_X2 _27623_ (.A(_22098_),
    .B(_22100_),
    .S(_04051_),
    .Z(_04262_));
 NOR3_X1 _27624_ (.A1(_04261_),
    .A2(_04262_),
    .A3(_04259_),
    .ZN(_04263_));
 NOR3_X1 _27625_ (.A1(_04234_),
    .A2(_04051_),
    .A3(_04229_),
    .ZN(_04264_));
 AOI21_X1 _27626_ (.A(_04079_),
    .B1(_04213_),
    .B2(_03974_),
    .ZN(_04265_));
 OAI21_X2 _27627_ (.A(_04203_),
    .B1(_03997_),
    .B2(_03982_),
    .ZN(_04266_));
 NOR2_X1 _27628_ (.A1(_04051_),
    .A2(_04226_),
    .ZN(_04267_));
 NAND2_X1 _27629_ (.A1(_04112_),
    .A2(_04104_),
    .ZN(_04268_));
 AOI221_X2 _27630_ (.A(_04264_),
    .B1(_04265_),
    .B2(_04266_),
    .C1(_04267_),
    .C2(_04268_),
    .ZN(_04269_));
 AOI211_X2 _27631_ (.A(_04259_),
    .B(_04263_),
    .C1(_04261_),
    .C2(_04269_),
    .ZN(_04270_));
 AOI211_X4 _27632_ (.A(_04226_),
    .B(_04212_),
    .C1(_04112_),
    .C2(_04104_),
    .ZN(_04271_));
 NOR2_X1 _27633_ (.A1(_04234_),
    .A2(_04229_),
    .ZN(_04272_));
 NAND2_X1 _27634_ (.A1(_04051_),
    .A2(_04209_),
    .ZN(_04273_));
 AOI21_X1 _27635_ (.A(_04273_),
    .B1(_04213_),
    .B2(_03974_),
    .ZN(_04274_));
 AOI221_X2 _27636_ (.A(_04271_),
    .B1(_04210_),
    .B2(_04272_),
    .C1(_04266_),
    .C2(_04274_),
    .ZN(_04275_));
 XNOR2_X2 _27637_ (.A(_04052_),
    .B(_04148_),
    .ZN(_04276_));
 NOR2_X2 _27638_ (.A1(_04152_),
    .A2(_04190_),
    .ZN(_04277_));
 NOR2_X2 _27639_ (.A1(_04276_),
    .A2(_04277_),
    .ZN(_04278_));
 AOI21_X4 _27640_ (.A(_04243_),
    .B1(_04275_),
    .B2(_04278_),
    .ZN(_04279_));
 NAND2_X1 _27641_ (.A1(_04240_),
    .A2(_04241_),
    .ZN(_04280_));
 OR4_X1 _27642_ (.A1(_04156_),
    .A2(_04204_),
    .A3(_04239_),
    .A4(_04280_),
    .ZN(_04281_));
 CLKBUF_X3 _27643_ (.A(_04281_),
    .Z(_04282_));
 OAI21_X2 _27644_ (.A(_04259_),
    .B1(_04279_),
    .B2(_04282_),
    .ZN(_04283_));
 NOR2_X2 _27645_ (.A1(_04252_),
    .A2(_04283_),
    .ZN(_04284_));
 BUF_X1 _27646_ (.A(_14162_),
    .Z(_04285_));
 INV_X2 _27647_ (.A(_04285_),
    .ZN(_04286_));
 BUF_X4 _27648_ (.A(_04286_),
    .Z(_14157_));
 OR2_X2 _27649_ (.A1(_04076_),
    .A2(_04113_),
    .ZN(_04287_));
 BUF_X4 _27650_ (.A(_04287_),
    .Z(_04288_));
 NOR2_X1 _27651_ (.A1(_04288_),
    .A2(_04269_),
    .ZN(_04289_));
 AOI21_X1 _27652_ (.A(_04289_),
    .B1(_04259_),
    .B2(_04191_),
    .ZN(_04290_));
 NOR2_X2 _27653_ (.A1(_14157_),
    .A2(_04290_),
    .ZN(_04291_));
 AOI21_X4 _27654_ (.A(_04270_),
    .B1(_04284_),
    .B2(_04291_),
    .ZN(_04292_));
 MUX2_X1 _27655_ (.A(_04249_),
    .B(_04247_),
    .S(_04257_),
    .Z(_04293_));
 CLKBUF_X3 _27656_ (.A(_04293_),
    .Z(_04294_));
 BUF_X4 _27657_ (.A(_04294_),
    .Z(_04295_));
 NAND3_X1 _27658_ (.A1(_04260_),
    .A2(_04182_),
    .A3(_04295_),
    .ZN(_04296_));
 OAI21_X1 _27659_ (.A(_04295_),
    .B1(_04262_),
    .B2(_04260_),
    .ZN(_04297_));
 NAND2_X1 _27660_ (.A1(_04140_),
    .A2(_04236_),
    .ZN(_04298_));
 AOI221_X2 _27661_ (.A(_04288_),
    .B1(_04139_),
    .B2(_04191_),
    .C1(_04207_),
    .C2(_04285_),
    .ZN(_04299_));
 XNOR2_X2 _27662_ (.A(_04257_),
    .B(_04138_),
    .ZN(_04300_));
 NOR4_X2 _27663_ (.A1(_04286_),
    .A2(_04288_),
    .A3(_04300_),
    .A4(_04269_),
    .ZN(_04301_));
 NAND2_X2 _27664_ (.A1(_04278_),
    .A2(_04275_),
    .ZN(_04302_));
 AOI22_X4 _27665_ (.A1(_04298_),
    .A2(_04299_),
    .B1(_04301_),
    .B2(_04302_),
    .ZN(_04303_));
 OAI211_X4 _27666_ (.A(_04259_),
    .B(_04253_),
    .C1(_04279_),
    .C2(_04282_),
    .ZN(_04304_));
 OAI21_X1 _27667_ (.A(_04297_),
    .B1(_04303_),
    .B2(_04304_),
    .ZN(_04305_));
 NAND2_X2 _27668_ (.A1(_04296_),
    .A2(_04305_),
    .ZN(_04306_));
 NOR2_X1 _27669_ (.A1(_04292_),
    .A2(_04306_),
    .ZN(_22110_));
 BUF_X4 _27670_ (.A(_03873_),
    .Z(_04307_));
 NOR4_X4 _27671_ (.A1(\g_reduce0[0].adder.x[11] ),
    .A2(\g_reduce0[0].adder.x[12] ),
    .A3(\g_reduce0[0].adder.x[14] ),
    .A4(_03871_),
    .ZN(_04308_));
 OR2_X1 _27672_ (.A1(_04308_),
    .A2(_03875_),
    .ZN(_04309_));
 CLKBUF_X3 _27673_ (.A(_04309_),
    .Z(_04310_));
 BUF_X4 _27674_ (.A(_04259_),
    .Z(_04311_));
 BUF_X4 _27675_ (.A(_04311_),
    .Z(_04312_));
 OR2_X1 _27676_ (.A1(_04294_),
    .A2(_04282_),
    .ZN(_04313_));
 OAI21_X4 _27677_ (.A(_04115_),
    .B1(_04279_),
    .B2(_04313_),
    .ZN(_04314_));
 NAND2_X1 _27678_ (.A1(_22105_),
    .A2(_22127_),
    .ZN(_04315_));
 OAI21_X1 _27679_ (.A(_04312_),
    .B1(_04314_),
    .B2(_04315_),
    .ZN(_04316_));
 NAND2_X1 _27680_ (.A1(_04306_),
    .A2(_04316_),
    .ZN(_04317_));
 MUX2_X1 _27681_ (.A(_04317_),
    .B(_04306_),
    .S(_04292_),
    .Z(_04318_));
 INV_X1 _27682_ (.A(_22112_),
    .ZN(_04319_));
 NOR2_X1 _27683_ (.A1(_04260_),
    .A2(_04115_),
    .ZN(_04320_));
 NAND2_X1 _27684_ (.A1(_04246_),
    .A2(_04276_),
    .ZN(_04321_));
 NAND2_X1 _27685_ (.A1(_04138_),
    .A2(_04276_),
    .ZN(_04322_));
 MUX2_X2 _27686_ (.A(_04321_),
    .B(_04322_),
    .S(_04117_),
    .Z(_04323_));
 NOR3_X2 _27687_ (.A1(_04288_),
    .A2(_04207_),
    .A3(_04323_),
    .ZN(_04324_));
 AOI211_X2 _27688_ (.A(_04287_),
    .B(_04182_),
    .C1(_04191_),
    .C2(_04139_),
    .ZN(_04325_));
 NAND2_X1 _27689_ (.A1(_04277_),
    .A2(_04262_),
    .ZN(_04326_));
 OAI21_X1 _27690_ (.A(_04286_),
    .B1(_04294_),
    .B2(_04326_),
    .ZN(_04327_));
 NOR3_X1 _27691_ (.A1(_04324_),
    .A2(_04325_),
    .A3(_04327_),
    .ZN(_04328_));
 NOR3_X2 _27692_ (.A1(_04288_),
    .A2(_04205_),
    .A3(_04323_),
    .ZN(_04329_));
 NAND2_X2 _27693_ (.A1(_04187_),
    .A2(_04186_),
    .ZN(_04330_));
 NAND3_X1 _27694_ (.A1(_04238_),
    .A2(_04161_),
    .A3(_04241_),
    .ZN(_04331_));
 NOR2_X1 _27695_ (.A1(_04169_),
    .A2(_04170_),
    .ZN(_04332_));
 AOI21_X1 _27696_ (.A(_04156_),
    .B1(_04161_),
    .B2(_04332_),
    .ZN(_04333_));
 NOR2_X1 _27697_ (.A1(_04152_),
    .A2(_04333_),
    .ZN(_04334_));
 NOR2_X2 _27698_ (.A1(_04276_),
    .A2(_04334_),
    .ZN(_04335_));
 NAND2_X1 _27699_ (.A1(_04331_),
    .A2(_04335_),
    .ZN(_04336_));
 AOI211_X2 _27700_ (.A(_04287_),
    .B(_04330_),
    .C1(_04336_),
    .C2(_04139_),
    .ZN(_04337_));
 NAND2_X1 _27701_ (.A1(_04181_),
    .A2(_04277_),
    .ZN(_04338_));
 NOR2_X2 _27702_ (.A1(_04294_),
    .A2(_04338_),
    .ZN(_04339_));
 NOR3_X2 _27703_ (.A1(_04329_),
    .A2(_04337_),
    .A3(_04339_),
    .ZN(_04340_));
 CLKBUF_X3 _27704_ (.A(_04285_),
    .Z(_04341_));
 AOI21_X2 _27705_ (.A(_04328_),
    .B1(_04340_),
    .B2(_04341_),
    .ZN(_04342_));
 MUX2_X1 _27706_ (.A(_04291_),
    .B(_04342_),
    .S(_22127_),
    .Z(_04343_));
 NOR3_X2 _27707_ (.A1(_04295_),
    .A2(_04279_),
    .A3(_04282_),
    .ZN(_04344_));
 NOR3_X1 _27708_ (.A1(_04161_),
    .A2(_04294_),
    .A3(_04335_),
    .ZN(_04345_));
 OAI21_X1 _27709_ (.A(_04140_),
    .B1(_04276_),
    .B2(_04238_),
    .ZN(_04346_));
 AND2_X1 _27710_ (.A1(_04114_),
    .A2(_04156_),
    .ZN(_04347_));
 AOI21_X2 _27711_ (.A(_04345_),
    .B1(_04346_),
    .B2(_04347_),
    .ZN(_04348_));
 OR3_X1 _27712_ (.A1(_14157_),
    .A2(_22127_),
    .A3(_04348_),
    .ZN(_04349_));
 NOR3_X1 _27713_ (.A1(_04138_),
    .A2(_04149_),
    .A3(_04241_),
    .ZN(_04350_));
 NOR3_X1 _27714_ (.A1(_04246_),
    .A2(_04149_),
    .A3(_04241_),
    .ZN(_04351_));
 MUX2_X1 _27715_ (.A(_04350_),
    .B(_04351_),
    .S(_04117_),
    .Z(_04352_));
 NOR3_X1 _27716_ (.A1(_04076_),
    .A2(_04113_),
    .A3(_04240_),
    .ZN(_04353_));
 NAND2_X1 _27717_ (.A1(_04246_),
    .A2(_04191_),
    .ZN(_04354_));
 NAND2_X1 _27718_ (.A1(_04138_),
    .A2(_04191_),
    .ZN(_04355_));
 MUX2_X1 _27719_ (.A(_04354_),
    .B(_04355_),
    .S(_04117_),
    .Z(_04356_));
 NOR3_X1 _27720_ (.A1(_04152_),
    .A2(_04241_),
    .A3(_04333_),
    .ZN(_04357_));
 AOI222_X2 _27721_ (.A1(_04115_),
    .A2(_04352_),
    .B1(_04353_),
    .B2(_04356_),
    .C1(_04357_),
    .C2(_04259_),
    .ZN(_04358_));
 NAND2_X1 _27722_ (.A1(_04140_),
    .A2(_04238_),
    .ZN(_04359_));
 NAND3_X1 _27723_ (.A1(_04115_),
    .A2(_04276_),
    .A3(_04359_),
    .ZN(_04360_));
 MUX2_X1 _27724_ (.A(_04358_),
    .B(_04360_),
    .S(_22127_),
    .Z(_04361_));
 OAI21_X1 _27725_ (.A(_04349_),
    .B1(_04361_),
    .B2(_04341_),
    .ZN(_04362_));
 AOI221_X2 _27726_ (.A(_04320_),
    .B1(_04343_),
    .B2(_04344_),
    .C1(_04362_),
    .C2(_04312_),
    .ZN(_04363_));
 INV_X1 _27727_ (.A(_04363_),
    .ZN(_04364_));
 CLKBUF_X3 _27728_ (.A(_04261_),
    .Z(_04365_));
 NOR2_X1 _27729_ (.A1(_04365_),
    .A2(_04115_),
    .ZN(_04366_));
 NOR2_X1 _27730_ (.A1(_04191_),
    .A2(_04236_),
    .ZN(_04367_));
 NOR2_X1 _27731_ (.A1(_04300_),
    .A2(_04335_),
    .ZN(_04368_));
 OAI33_X1 _27732_ (.A1(_04330_),
    .A2(_04367_),
    .A3(_04295_),
    .B1(_04368_),
    .B2(_04288_),
    .B3(_04241_),
    .ZN(_04369_));
 NOR2_X1 _27733_ (.A1(_04341_),
    .A2(_04253_),
    .ZN(_04370_));
 MUX2_X1 _27734_ (.A(_04276_),
    .B(_04156_),
    .S(_04286_),
    .Z(_04371_));
 NOR2_X1 _27735_ (.A1(_04341_),
    .A2(_04238_),
    .ZN(_04372_));
 AOI22_X1 _27736_ (.A1(_04140_),
    .A2(_04371_),
    .B1(_04372_),
    .B2(_04323_),
    .ZN(_04373_));
 MUX2_X1 _27737_ (.A(_04240_),
    .B(_04161_),
    .S(_04237_),
    .Z(_04374_));
 NAND2_X1 _27738_ (.A1(_04341_),
    .A2(_04252_),
    .ZN(_04375_));
 OAI22_X1 _27739_ (.A1(_04252_),
    .A2(_04373_),
    .B1(_04374_),
    .B2(_04375_),
    .ZN(_04376_));
 AOI221_X2 _27740_ (.A(_04314_),
    .B1(_04369_),
    .B2(_04370_),
    .C1(_04376_),
    .C2(_04115_),
    .ZN(_04377_));
 NOR3_X1 _27741_ (.A1(_04288_),
    .A2(_04191_),
    .A3(_04207_),
    .ZN(_04378_));
 NOR2_X1 _27742_ (.A1(_04191_),
    .A2(_04209_),
    .ZN(_04379_));
 OAI33_X1 _27743_ (.A1(_04288_),
    .A2(_04140_),
    .A3(_04207_),
    .B1(_04269_),
    .B2(_04294_),
    .B3(_04379_),
    .ZN(_04380_));
 NOR2_X2 _27744_ (.A1(_04378_),
    .A2(_04380_),
    .ZN(_04381_));
 NAND2_X2 _27745_ (.A1(_14157_),
    .A2(_04253_),
    .ZN(_04382_));
 NAND2_X1 _27746_ (.A1(_04341_),
    .A2(_04253_),
    .ZN(_04383_));
 NOR3_X1 _27747_ (.A1(_04287_),
    .A2(_04182_),
    .A3(_04323_),
    .ZN(_04384_));
 NOR2_X1 _27748_ (.A1(_04182_),
    .A2(_04294_),
    .ZN(_04385_));
 OR2_X1 _27749_ (.A1(_04277_),
    .A2(_04236_),
    .ZN(_04386_));
 OAI21_X1 _27750_ (.A(_04335_),
    .B1(_04331_),
    .B2(_04330_),
    .ZN(_04387_));
 NAND2_X1 _27751_ (.A1(_04139_),
    .A2(_04387_),
    .ZN(_04388_));
 NOR2_X1 _27752_ (.A1(_04287_),
    .A2(_04205_),
    .ZN(_04389_));
 AOI221_X2 _27753_ (.A(_04384_),
    .B1(_04385_),
    .B2(_04386_),
    .C1(_04388_),
    .C2(_04389_),
    .ZN(_04390_));
 OAI22_X4 _27754_ (.A1(_04381_),
    .A2(_04382_),
    .B1(_04383_),
    .B2(_04390_),
    .ZN(_04391_));
 AOI21_X1 _27755_ (.A(_04391_),
    .B1(_04252_),
    .B2(_22105_),
    .ZN(_04392_));
 AOI21_X1 _27756_ (.A(_04377_),
    .B1(_04392_),
    .B2(_04314_),
    .ZN(_04393_));
 AOI221_X2 _27757_ (.A(_04366_),
    .B1(_04393_),
    .B2(_04311_),
    .C1(_04365_),
    .C2(_04300_),
    .ZN(_04394_));
 OAI211_X2 _27758_ (.A(_04259_),
    .B(_04252_),
    .C1(_04279_),
    .C2(_04282_),
    .ZN(_04395_));
 AND2_X1 _27759_ (.A1(_04341_),
    .A2(_04358_),
    .ZN(_04396_));
 NOR4_X2 _27760_ (.A1(_04341_),
    .A2(_04329_),
    .A3(_04337_),
    .A4(_04339_),
    .ZN(_04397_));
 NOR3_X1 _27761_ (.A1(_04395_),
    .A2(_04396_),
    .A3(_04397_),
    .ZN(_04398_));
 MUX2_X1 _27762_ (.A(_04360_),
    .B(_04348_),
    .S(_14157_),
    .Z(_04399_));
 NAND2_X1 _27763_ (.A1(_04285_),
    .A2(_04182_),
    .ZN(_04400_));
 NOR2_X1 _27764_ (.A1(_04276_),
    .A2(_04400_),
    .ZN(_04401_));
 NOR3_X1 _27765_ (.A1(_04286_),
    .A2(_04300_),
    .A3(_04262_),
    .ZN(_04402_));
 MUX2_X1 _27766_ (.A(_04401_),
    .B(_04402_),
    .S(_04386_),
    .Z(_04403_));
 NAND3_X1 _27767_ (.A1(_04286_),
    .A2(_04269_),
    .A3(_04356_),
    .ZN(_04404_));
 OR2_X1 _27768_ (.A1(_04140_),
    .A2(_04400_),
    .ZN(_04405_));
 NAND4_X1 _27769_ (.A1(_04285_),
    .A2(_04140_),
    .A3(_04276_),
    .A4(_04207_),
    .ZN(_04406_));
 NAND4_X1 _27770_ (.A1(_04115_),
    .A2(_04404_),
    .A3(_04405_),
    .A4(_04406_),
    .ZN(_04407_));
 OR2_X1 _27771_ (.A1(_04403_),
    .A2(_04407_),
    .ZN(_04408_));
 XNOR2_X1 _27772_ (.A(_22107_),
    .B(_04245_),
    .ZN(_04409_));
 NAND2_X1 _27773_ (.A1(_04344_),
    .A2(_04409_),
    .ZN(_04410_));
 MUX2_X1 _27774_ (.A(_04140_),
    .B(_04149_),
    .S(_04365_),
    .Z(_04411_));
 OAI222_X2 _27775_ (.A1(_04304_),
    .A2(_04399_),
    .B1(_04408_),
    .B2(_04410_),
    .C1(_04411_),
    .C2(_04311_),
    .ZN(_04412_));
 OR2_X1 _27776_ (.A1(_04398_),
    .A2(_04412_),
    .ZN(_04413_));
 MUX2_X1 _27777_ (.A(_04152_),
    .B(_04156_),
    .S(_04365_),
    .Z(_04414_));
 NOR2_X1 _27778_ (.A1(_04311_),
    .A2(_04414_),
    .ZN(_04415_));
 NOR2_X1 _27779_ (.A1(_04358_),
    .A2(_04382_),
    .ZN(_04416_));
 NAND2_X1 _27780_ (.A1(_04252_),
    .A2(_04340_),
    .ZN(_04417_));
 AOI21_X1 _27781_ (.A(_14157_),
    .B1(_04253_),
    .B2(_04348_),
    .ZN(_04418_));
 NOR2_X1 _27782_ (.A1(_04295_),
    .A2(_04326_),
    .ZN(_04419_));
 OR3_X1 _27783_ (.A1(_04324_),
    .A2(_04325_),
    .A3(_04419_),
    .ZN(_04420_));
 AOI221_X2 _27784_ (.A(_04416_),
    .B1(_04417_),
    .B2(_04418_),
    .C1(_04370_),
    .C2(_04420_),
    .ZN(_04421_));
 NOR2_X4 _27785_ (.A1(_04295_),
    .A2(_04314_),
    .ZN(_04422_));
 INV_X1 _27786_ (.A(_04314_),
    .ZN(_22131_));
 AOI21_X1 _27787_ (.A(_22131_),
    .B1(_04291_),
    .B2(_22127_),
    .ZN(_04423_));
 AOI221_X2 _27788_ (.A(_04415_),
    .B1(_04421_),
    .B2(_04422_),
    .C1(_04423_),
    .C2(_04311_),
    .ZN(_04424_));
 NOR2_X1 _27789_ (.A1(_22127_),
    .A2(_04390_),
    .ZN(_04425_));
 NAND2_X1 _27790_ (.A1(_04115_),
    .A2(_22127_),
    .ZN(_04426_));
 OAI21_X1 _27791_ (.A(_14157_),
    .B1(_04374_),
    .B2(_04426_),
    .ZN(_04427_));
 AOI22_X1 _27792_ (.A1(_04140_),
    .A2(_04156_),
    .B1(_04323_),
    .B2(_04152_),
    .ZN(_04428_));
 NOR2_X1 _27793_ (.A1(_04288_),
    .A2(_04428_),
    .ZN(_04429_));
 MUX2_X1 _27794_ (.A(_04369_),
    .B(_04429_),
    .S(_22127_),
    .Z(_04430_));
 OAI221_X2 _27795_ (.A(_04422_),
    .B1(_04425_),
    .B2(_04427_),
    .C1(_04430_),
    .C2(_14157_),
    .ZN(_04431_));
 MUX2_X1 _27796_ (.A(_04149_),
    .B(_04238_),
    .S(_04365_),
    .Z(_04432_));
 OAI221_X2 _27797_ (.A(_04431_),
    .B1(_04410_),
    .B2(_04303_),
    .C1(_04311_),
    .C2(_04432_),
    .ZN(_04433_));
 NAND3_X1 _27798_ (.A1(_04413_),
    .A2(_04424_),
    .A3(_04433_),
    .ZN(_04434_));
 NAND2_X1 _27799_ (.A1(_22105_),
    .A2(_04252_),
    .ZN(_04435_));
 MUX2_X1 _27800_ (.A(_04330_),
    .B(_04205_),
    .S(_04261_),
    .Z(_04436_));
 OAI22_X2 _27801_ (.A1(_04283_),
    .A2(_04435_),
    .B1(_04436_),
    .B2(_04311_),
    .ZN(_04437_));
 AOI21_X4 _27802_ (.A(_04437_),
    .B1(_04391_),
    .B2(_04422_),
    .ZN(_04438_));
 NOR3_X1 _27803_ (.A1(_04304_),
    .A2(_04403_),
    .A3(_04407_),
    .ZN(_04439_));
 MUX2_X1 _27804_ (.A(_04205_),
    .B(_04182_),
    .S(_04261_),
    .Z(_04440_));
 NOR2_X1 _27805_ (.A1(_04311_),
    .A2(_04440_),
    .ZN(_04441_));
 NOR2_X2 _27806_ (.A1(_04439_),
    .A2(_04441_),
    .ZN(_04442_));
 NOR4_X4 _27807_ (.A1(_04292_),
    .A2(_04306_),
    .A3(_04438_),
    .A4(_04442_),
    .ZN(_04443_));
 NOR3_X2 _27808_ (.A1(_04304_),
    .A2(_04396_),
    .A3(_04397_),
    .ZN(_04444_));
 MUX2_X1 _27809_ (.A(_04161_),
    .B(_04240_),
    .S(_04261_),
    .Z(_04445_));
 NOR2_X1 _27810_ (.A1(_04257_),
    .A2(_04249_),
    .ZN(_04446_));
 NOR2_X1 _27811_ (.A1(_04117_),
    .A2(_04247_),
    .ZN(_04447_));
 OAI33_X1 _27812_ (.A1(_04395_),
    .A2(_04403_),
    .A3(_04407_),
    .B1(_04445_),
    .B2(_04446_),
    .B3(_04447_),
    .ZN(_04448_));
 MUX2_X1 _27813_ (.A(_04176_),
    .B(_04242_),
    .S(_04261_),
    .Z(_04449_));
 NAND2_X1 _27814_ (.A1(_04295_),
    .A2(_04449_),
    .ZN(_04450_));
 AOI21_X1 _27815_ (.A(_04387_),
    .B1(_04289_),
    .B2(_04282_),
    .ZN(_04451_));
 NAND3_X1 _27816_ (.A1(_04341_),
    .A2(_04259_),
    .A3(_04252_),
    .ZN(_04452_));
 OAI21_X1 _27817_ (.A(_04285_),
    .B1(_04295_),
    .B2(_04338_),
    .ZN(_04453_));
 OAI33_X1 _27818_ (.A1(_04329_),
    .A2(_04337_),
    .A3(_04453_),
    .B1(_04324_),
    .B2(_04325_),
    .B3(_04327_),
    .ZN(_04454_));
 OAI221_X2 _27819_ (.A(_04450_),
    .B1(_04451_),
    .B2(_04452_),
    .C1(_04454_),
    .C2(_04304_),
    .ZN(_04455_));
 AOI22_X2 _27820_ (.A1(_04342_),
    .A2(_04444_),
    .B1(_04448_),
    .B2(_04455_),
    .ZN(_04456_));
 MUX2_X1 _27821_ (.A(_04240_),
    .B(_04241_),
    .S(_04261_),
    .Z(_04457_));
 OAI22_X2 _27822_ (.A1(_04303_),
    .A2(_04395_),
    .B1(_04457_),
    .B2(_04311_),
    .ZN(_04458_));
 OR2_X1 _27823_ (.A1(_04300_),
    .A2(_04335_),
    .ZN(_04459_));
 NOR2_X1 _27824_ (.A1(_04288_),
    .A2(_04241_),
    .ZN(_04460_));
 NOR2_X1 _27825_ (.A1(_04330_),
    .A2(_04294_),
    .ZN(_04461_));
 AOI221_X2 _27826_ (.A(_04286_),
    .B1(_04459_),
    .B2(_04460_),
    .C1(_04461_),
    .C2(_04302_),
    .ZN(_04462_));
 AOI21_X2 _27827_ (.A(_04462_),
    .B1(_04390_),
    .B2(_14157_),
    .ZN(_04463_));
 AOI21_X4 _27828_ (.A(_04458_),
    .B1(_04463_),
    .B2(_04284_),
    .ZN(_04464_));
 MUX2_X1 _27829_ (.A(_04156_),
    .B(_04204_),
    .S(_04365_),
    .Z(_04465_));
 NAND2_X1 _27830_ (.A1(_04295_),
    .A2(_04465_),
    .ZN(_04466_));
 AOI21_X1 _27831_ (.A(_04295_),
    .B1(_04314_),
    .B2(_04315_),
    .ZN(_04467_));
 AOI22_X1 _27832_ (.A1(_04459_),
    .A2(_04460_),
    .B1(_04461_),
    .B2(_04302_),
    .ZN(_04468_));
 NAND2_X1 _27833_ (.A1(_14157_),
    .A2(_04252_),
    .ZN(_04469_));
 OAI221_X1 _27834_ (.A(_22131_),
    .B1(_04382_),
    .B2(_04468_),
    .C1(_04469_),
    .C2(_04381_),
    .ZN(_04470_));
 NAND3_X1 _27835_ (.A1(_04341_),
    .A2(_04115_),
    .A3(_22127_),
    .ZN(_04471_));
 OAI22_X1 _27836_ (.A1(_04390_),
    .A2(_04375_),
    .B1(_04471_),
    .B2(_04374_),
    .ZN(_04472_));
 OAI21_X1 _27837_ (.A(_04467_),
    .B1(_04470_),
    .B2(_04472_),
    .ZN(_04473_));
 AOI211_X2 _27838_ (.A(_04456_),
    .B(_04464_),
    .C1(_04466_),
    .C2(_04473_),
    .ZN(_04474_));
 NAND2_X2 _27839_ (.A1(_04443_),
    .A2(_04474_),
    .ZN(_04475_));
 OR3_X1 _27840_ (.A1(_04394_),
    .A2(_04434_),
    .A3(_04475_),
    .ZN(_04476_));
 XNOR2_X1 _27841_ (.A(_04364_),
    .B(_04476_),
    .ZN(_22115_));
 MUX2_X1 _27842_ (.A(_04318_),
    .B(_04319_),
    .S(_22115_),
    .Z(_04477_));
 NAND2_X4 _27843_ (.A1(_03873_),
    .A2(_03875_),
    .ZN(_04478_));
 OAI222_X2 _27844_ (.A1(_03899_),
    .A2(_04307_),
    .B1(_04310_),
    .B2(_04477_),
    .C1(_04478_),
    .C2(_03922_),
    .ZN(_00128_));
 XNOR2_X1 _27845_ (.A(_22111_),
    .B(_04438_),
    .ZN(_04479_));
 NOR2_X1 _27846_ (.A1(_04310_),
    .A2(_04479_),
    .ZN(_04480_));
 AND2_X1 _27847_ (.A1(_22115_),
    .A2(_04480_),
    .ZN(_04481_));
 NOR3_X1 _27848_ (.A1(_22112_),
    .A2(_04310_),
    .A3(_22115_),
    .ZN(_04482_));
 OAI22_X2 _27849_ (.A1(\g_reduce0[2].adder.x[1] ),
    .A2(_03873_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[1] ),
    .ZN(_04483_));
 NOR3_X1 _27850_ (.A1(_04481_),
    .A2(_04482_),
    .A3(_04483_),
    .ZN(_00135_));
 OAI22_X2 _27851_ (.A1(\g_reduce0[2].adder.x[2] ),
    .A2(_04307_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[2] ),
    .ZN(_04484_));
 INV_X1 _27852_ (.A(_04455_),
    .ZN(_04485_));
 XNOR2_X1 _27853_ (.A(_04443_),
    .B(_04485_),
    .ZN(_04486_));
 NOR2_X1 _27854_ (.A1(_04310_),
    .A2(_04486_),
    .ZN(_04487_));
 MUX2_X1 _27855_ (.A(_04480_),
    .B(_04487_),
    .S(_22115_),
    .Z(_04488_));
 NOR2_X1 _27856_ (.A1(_04484_),
    .A2(_04488_),
    .ZN(_00136_));
 OAI22_X2 _27857_ (.A1(\g_reduce0[2].adder.x[3] ),
    .A2(_04307_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[3] ),
    .ZN(_04489_));
 INV_X1 _27858_ (.A(_22111_),
    .ZN(_04490_));
 NOR2_X2 _27859_ (.A1(_04490_),
    .A2(_04438_),
    .ZN(_04491_));
 NAND2_X1 _27860_ (.A1(_04455_),
    .A2(_04491_),
    .ZN(_04492_));
 XOR2_X1 _27861_ (.A(_04464_),
    .B(_04492_),
    .Z(_04493_));
 NOR2_X1 _27862_ (.A1(_04310_),
    .A2(_04493_),
    .ZN(_04494_));
 MUX2_X1 _27863_ (.A(_04487_),
    .B(_04494_),
    .S(_22115_),
    .Z(_04495_));
 NOR2_X1 _27864_ (.A1(_04489_),
    .A2(_04495_),
    .ZN(_00137_));
 OAI22_X2 _27865_ (.A1(\g_reduce0[2].adder.x[4] ),
    .A2(_04307_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[4] ),
    .ZN(_04496_));
 NOR2_X1 _27866_ (.A1(_04456_),
    .A2(_04464_),
    .ZN(_04497_));
 NAND2_X1 _27867_ (.A1(_04443_),
    .A2(_04497_),
    .ZN(_04498_));
 NOR2_X1 _27868_ (.A1(_04444_),
    .A2(_04448_),
    .ZN(_04499_));
 OR2_X1 _27869_ (.A1(_04485_),
    .A2(_04464_),
    .ZN(_04500_));
 INV_X1 _27870_ (.A(_04443_),
    .ZN(_04501_));
 OAI21_X1 _27871_ (.A(_04499_),
    .B1(_04500_),
    .B2(_04501_),
    .ZN(_04502_));
 AOI21_X1 _27872_ (.A(_04309_),
    .B1(_04498_),
    .B2(_04502_),
    .ZN(_04503_));
 MUX2_X1 _27873_ (.A(_04494_),
    .B(_04503_),
    .S(_22115_),
    .Z(_04504_));
 NOR2_X1 _27874_ (.A1(_04496_),
    .A2(_04504_),
    .ZN(_00138_));
 AND2_X1 _27875_ (.A1(_04466_),
    .A2(_04473_),
    .ZN(_04505_));
 AND2_X1 _27876_ (.A1(_04497_),
    .A2(_04491_),
    .ZN(_04506_));
 XNOR2_X1 _27877_ (.A(_04505_),
    .B(_04506_),
    .ZN(_04507_));
 NOR2_X1 _27878_ (.A1(_04310_),
    .A2(_04507_),
    .ZN(_04508_));
 MUX2_X1 _27879_ (.A(_04503_),
    .B(_04508_),
    .S(_22115_),
    .Z(_04509_));
 OAI22_X2 _27880_ (.A1(\g_reduce0[2].adder.x[5] ),
    .A2(_04307_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[5] ),
    .ZN(_04510_));
 NOR2_X1 _27881_ (.A1(_04509_),
    .A2(_04510_),
    .ZN(_00139_));
 OAI22_X2 _27882_ (.A1(\g_reduce0[2].adder.x[6] ),
    .A2(_03873_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[6] ),
    .ZN(_04511_));
 AND2_X1 _27883_ (.A1(_04476_),
    .A2(_04507_),
    .ZN(_04512_));
 AOI21_X1 _27884_ (.A(_04310_),
    .B1(_04363_),
    .B2(_04512_),
    .ZN(_04513_));
 XNOR2_X2 _27885_ (.A(_04424_),
    .B(_04475_),
    .ZN(_04514_));
 OR2_X1 _27886_ (.A1(_04394_),
    .A2(_04434_),
    .ZN(_04515_));
 NOR4_X1 _27887_ (.A1(_04515_),
    .A2(_04505_),
    .A3(_04498_),
    .A4(_04506_),
    .ZN(_04516_));
 OAI21_X1 _27888_ (.A(_04364_),
    .B1(_04514_),
    .B2(_04516_),
    .ZN(_04517_));
 AOI21_X1 _27889_ (.A(_04511_),
    .B1(_04513_),
    .B2(_04517_),
    .ZN(_00140_));
 AND2_X1 _27890_ (.A1(_04474_),
    .A2(_04491_),
    .ZN(_04518_));
 NAND2_X1 _27891_ (.A1(_04424_),
    .A2(_04518_),
    .ZN(_04519_));
 XNOR2_X1 _27892_ (.A(_04433_),
    .B(_04519_),
    .ZN(_04520_));
 AOI221_X2 _27893_ (.A(_04309_),
    .B1(_04363_),
    .B2(_04514_),
    .C1(_04520_),
    .C2(_22115_),
    .ZN(_04521_));
 OAI22_X2 _27894_ (.A1(\g_reduce0[2].adder.x[7] ),
    .A2(_04307_),
    .B1(_04478_),
    .B2(\g_reduce0[0].adder.x[7] ),
    .ZN(_04522_));
 NOR2_X1 _27895_ (.A1(_04521_),
    .A2(_04522_),
    .ZN(_00141_));
 AND2_X1 _27896_ (.A1(_03873_),
    .A2(_03875_),
    .ZN(_04523_));
 AOI22_X2 _27897_ (.A1(\g_reduce0[2].adder.x[8] ),
    .A2(_04308_),
    .B1(_04523_),
    .B2(\g_reduce0[0].adder.x[8] ),
    .ZN(_04524_));
 XOR2_X1 _27898_ (.A(_04433_),
    .B(_04519_),
    .Z(_04525_));
 NAND2_X1 _27899_ (.A1(_04424_),
    .A2(_04433_),
    .ZN(_04526_));
 NOR2_X1 _27900_ (.A1(_04526_),
    .A2(_04475_),
    .ZN(_04527_));
 XNOR2_X1 _27901_ (.A(_04413_),
    .B(_04527_),
    .ZN(_04528_));
 MUX2_X1 _27902_ (.A(_04525_),
    .B(_04528_),
    .S(_22115_),
    .Z(_04529_));
 OAI21_X1 _27903_ (.A(_04524_),
    .B1(_04529_),
    .B2(_04310_),
    .ZN(_00142_));
 NAND2_X1 _27904_ (.A1(_04474_),
    .A2(_04491_),
    .ZN(_04530_));
 OAI21_X1 _27905_ (.A(_04394_),
    .B1(_04434_),
    .B2(_04530_),
    .ZN(_04531_));
 OAI21_X1 _27906_ (.A(_04474_),
    .B1(_04491_),
    .B2(_04443_),
    .ZN(_04532_));
 OAI21_X1 _27907_ (.A(_04531_),
    .B1(_04532_),
    .B2(_04515_),
    .ZN(_04533_));
 NOR3_X1 _27908_ (.A1(_04310_),
    .A2(_04363_),
    .A3(_04533_),
    .ZN(_04534_));
 NOR2_X1 _27909_ (.A1(_04413_),
    .A2(_04527_),
    .ZN(_04535_));
 OAI21_X1 _27910_ (.A(_04413_),
    .B1(_04518_),
    .B2(_04394_),
    .ZN(_04536_));
 NOR3_X1 _27911_ (.A1(_04526_),
    .A2(_04475_),
    .A3(_04536_),
    .ZN(_04537_));
 NOR4_X1 _27912_ (.A1(_04310_),
    .A2(_04364_),
    .A3(_04535_),
    .A4(_04537_),
    .ZN(_04538_));
 AOI22_X2 _27913_ (.A1(\g_reduce0[2].adder.x[9] ),
    .A2(_04308_),
    .B1(_04523_),
    .B2(\g_reduce0[0].adder.x[9] ),
    .ZN(_04539_));
 INV_X1 _27914_ (.A(_04539_),
    .ZN(_04540_));
 OR3_X1 _27915_ (.A1(_04534_),
    .A2(_04538_),
    .A3(_04540_),
    .ZN(_00143_));
 INV_X1 _27916_ (.A(_22119_),
    .ZN(_22113_));
 MUX2_X1 _27917_ (.A(_22118_),
    .B(\g_reduce0[0].adder.x[10] ),
    .S(_03875_),
    .Z(_04541_));
 MUX2_X1 _27918_ (.A(\g_reduce0[2].adder.x[10] ),
    .B(_04541_),
    .S(_04307_),
    .Z(_00129_));
 MUX2_X1 _27919_ (.A(_22126_),
    .B(\g_reduce0[0].adder.x[11] ),
    .S(_03875_),
    .Z(_04542_));
 MUX2_X1 _27920_ (.A(\g_reduce0[2].adder.x[11] ),
    .B(_04542_),
    .S(_04307_),
    .Z(_00130_));
 MUX2_X2 _27921_ (.A(_21994_),
    .B(_00570_),
    .S(_03931_),
    .Z(_04543_));
 NAND2_X1 _27922_ (.A1(_04260_),
    .A2(_22120_),
    .ZN(_04544_));
 XOR2_X1 _27923_ (.A(_04543_),
    .B(_04544_),
    .Z(_04545_));
 XNOR2_X1 _27924_ (.A(_14160_),
    .B(_22130_),
    .ZN(_04546_));
 MUX2_X1 _27925_ (.A(_04545_),
    .B(_04546_),
    .S(_04311_),
    .Z(_04547_));
 XOR2_X1 _27926_ (.A(_22125_),
    .B(_04547_),
    .Z(_04548_));
 MUX2_X1 _27927_ (.A(_04548_),
    .B(\g_reduce0[0].adder.x[12] ),
    .S(_03875_),
    .Z(_04549_));
 MUX2_X1 _27928_ (.A(\g_reduce0[2].adder.x[12] ),
    .B(_04549_),
    .S(_04307_),
    .Z(_00131_));
 MUX2_X1 _27929_ (.A(_21991_),
    .B(_00573_),
    .S(_03935_),
    .Z(_04550_));
 NOR4_X1 _27930_ (.A1(_04365_),
    .A2(_22113_),
    .A3(_14159_),
    .A4(_04543_),
    .ZN(_04551_));
 XNOR2_X1 _27931_ (.A(_04550_),
    .B(_04551_),
    .ZN(_04552_));
 INV_X1 _27932_ (.A(_22129_),
    .ZN(_04553_));
 INV_X1 _27933_ (.A(_14158_),
    .ZN(_04554_));
 AOI21_X1 _27934_ (.A(_22122_),
    .B1(_22123_),
    .B2(_04554_),
    .ZN(_04555_));
 INV_X1 _27935_ (.A(_22130_),
    .ZN(_04556_));
 OAI21_X1 _27936_ (.A(_04553_),
    .B1(_04555_),
    .B2(_04556_),
    .ZN(_04557_));
 XOR2_X1 _27937_ (.A(_22134_),
    .B(_04557_),
    .Z(_04558_));
 MUX2_X1 _27938_ (.A(_04552_),
    .B(_04558_),
    .S(_04312_),
    .Z(_04559_));
 NOR2_X1 _27939_ (.A1(_04365_),
    .A2(_22121_),
    .ZN(_04560_));
 AOI21_X1 _27940_ (.A(_04560_),
    .B1(_14159_),
    .B2(_04365_),
    .ZN(_04561_));
 NOR2_X1 _27941_ (.A1(_04312_),
    .A2(_04561_),
    .ZN(_04562_));
 AOI21_X2 _27942_ (.A(_04562_),
    .B1(_04312_),
    .B2(_14161_),
    .ZN(_22124_));
 NAND3_X1 _27943_ (.A1(_22117_),
    .A2(_04547_),
    .A3(_22124_),
    .ZN(_04563_));
 XNOR2_X1 _27944_ (.A(_04559_),
    .B(_04563_),
    .ZN(_04564_));
 MUX2_X1 _27945_ (.A(_04564_),
    .B(\g_reduce0[0].adder.x[13] ),
    .S(_03875_),
    .Z(_04565_));
 MUX2_X1 _27946_ (.A(\g_reduce0[2].adder.x[13] ),
    .B(_04565_),
    .S(_03873_),
    .Z(_00132_));
 BUF_X4 _27947_ (.A(_03935_),
    .Z(_04566_));
 NOR4_X1 _27948_ (.A1(_04312_),
    .A2(_04543_),
    .A3(_04544_),
    .A4(_04550_),
    .ZN(_04567_));
 OAI21_X1 _27949_ (.A(_04553_),
    .B1(_04556_),
    .B2(_14160_),
    .ZN(_04568_));
 AOI21_X1 _27950_ (.A(_22133_),
    .B1(_04568_),
    .B2(_22134_),
    .ZN(_04569_));
 AOI21_X1 _27951_ (.A(_04567_),
    .B1(_04569_),
    .B2(_04312_),
    .ZN(_04570_));
 NAND3_X1 _27952_ (.A1(_22125_),
    .A2(_04547_),
    .A3(_04559_),
    .ZN(_04571_));
 XOR2_X2 _27953_ (.A(_04570_),
    .B(_04571_),
    .Z(_04572_));
 AND3_X1 _27954_ (.A1(\g_reduce0[2].adder.x[14] ),
    .A2(_04566_),
    .A3(_04572_),
    .ZN(_04573_));
 NOR2_X1 _27955_ (.A1(_04566_),
    .A2(_04572_),
    .ZN(_04574_));
 NOR3_X1 _27956_ (.A1(_03875_),
    .A2(_04573_),
    .A3(_04574_),
    .ZN(_04575_));
 NOR3_X1 _27957_ (.A1(\g_reduce0[0].adder.x[14] ),
    .A2(_04308_),
    .A3(_04575_),
    .ZN(_04576_));
 OR2_X1 _27958_ (.A1(\g_reduce0[2].adder.x[14] ),
    .A2(_03908_),
    .ZN(_04577_));
 NAND2_X1 _27959_ (.A1(\g_reduce0[0].adder.x[14] ),
    .A2(_04577_),
    .ZN(_04578_));
 MUX2_X1 _27960_ (.A(_04577_),
    .B(_04578_),
    .S(_04572_),
    .Z(_04579_));
 OAI22_X1 _27961_ (.A1(\g_reduce0[2].adder.x[14] ),
    .A2(_04307_),
    .B1(_03875_),
    .B2(_04579_),
    .ZN(_04580_));
 NOR2_X1 _27962_ (.A1(_04576_),
    .A2(_04580_),
    .ZN(_00133_));
 BUF_X2 _27963_ (.A(\g_reduce0[4].adder.x[11] ),
    .Z(_04581_));
 BUF_X2 _27964_ (.A(\g_reduce0[4].adder.x[12] ),
    .Z(_04582_));
 BUF_X2 _27965_ (.A(\g_reduce0[4].adder.x[14] ),
    .Z(_04583_));
 OR2_X2 _27966_ (.A1(\g_reduce0[4].adder.x[10] ),
    .A2(\g_reduce0[4].adder.x[13] ),
    .ZN(_04584_));
 OR4_X4 _27967_ (.A1(_04581_),
    .A2(_04582_),
    .A3(_04583_),
    .A4(_04584_),
    .ZN(_04585_));
 INV_X1 _27968_ (.A(\g_reduce0[6].adder.x[14] ),
    .ZN(_04586_));
 NOR4_X1 _27969_ (.A1(\g_reduce0[6].adder.x[11] ),
    .A2(\g_reduce0[6].adder.x[10] ),
    .A3(\g_reduce0[6].adder.x[13] ),
    .A4(\g_reduce0[6].adder.x[12] ),
    .ZN(_04587_));
 AND2_X1 _27970_ (.A1(_04586_),
    .A2(_04587_),
    .ZN(_04588_));
 BUF_X4 _27971_ (.A(_04588_),
    .Z(_04589_));
 INV_X1 _27972_ (.A(_22181_),
    .ZN(_04590_));
 BUF_X2 _27973_ (.A(_22137_),
    .Z(_04591_));
 AOI21_X2 _27974_ (.A(_22136_),
    .B1(_22139_),
    .B2(_04591_),
    .ZN(_04592_));
 BUF_X2 _27975_ (.A(_22182_),
    .Z(_04593_));
 INV_X1 _27976_ (.A(_04593_),
    .ZN(_04594_));
 OAI21_X2 _27977_ (.A(_04590_),
    .B1(_04592_),
    .B2(_04594_),
    .ZN(_04595_));
 INV_X1 _27978_ (.A(_22142_),
    .ZN(_04596_));
 BUF_X1 _27979_ (.A(_22143_),
    .Z(_04597_));
 INV_X1 _27980_ (.A(_04597_),
    .ZN(_04598_));
 OAI21_X2 _27981_ (.A(_04596_),
    .B1(_22175_),
    .B2(_04598_),
    .ZN(_04599_));
 CLKBUF_X3 _27982_ (.A(_22140_),
    .Z(_04600_));
 AND2_X1 _27983_ (.A1(_04591_),
    .A2(_04600_),
    .ZN(_04601_));
 AND2_X1 _27984_ (.A1(_04593_),
    .A2(_04601_),
    .ZN(_04602_));
 AOI21_X4 _27985_ (.A(_04595_),
    .B1(_04599_),
    .B2(_04602_),
    .ZN(_04603_));
 BUF_X2 _27986_ (.A(_22176_),
    .Z(_04604_));
 INV_X1 _27987_ (.A(_04604_),
    .ZN(_04605_));
 NAND3_X2 _27988_ (.A1(_04593_),
    .A2(_04591_),
    .A3(_04600_),
    .ZN(_04606_));
 NOR3_X4 _27989_ (.A1(_04605_),
    .A2(_04598_),
    .A3(_04606_),
    .ZN(_04607_));
 AOI21_X1 _27990_ (.A(_22145_),
    .B1(_22148_),
    .B2(_22146_),
    .ZN(_04608_));
 AOI21_X1 _27991_ (.A(_22151_),
    .B1(_22152_),
    .B2(_22154_),
    .ZN(_04609_));
 NAND2_X1 _27992_ (.A1(_22146_),
    .A2(_22149_),
    .ZN(_04610_));
 OAI21_X1 _27993_ (.A(_04608_),
    .B1(_04609_),
    .B2(_04610_),
    .ZN(_04611_));
 INV_X1 _27994_ (.A(_22169_),
    .ZN(_04612_));
 INV_X1 _27995_ (.A(_22170_),
    .ZN(_04613_));
 OAI21_X1 _27996_ (.A(_04612_),
    .B1(_22172_),
    .B2(_04613_),
    .ZN(_04614_));
 AND4_X1 _27997_ (.A1(_22146_),
    .A2(_22149_),
    .A3(_22152_),
    .A4(_22155_),
    .ZN(_04615_));
 AND3_X1 _27998_ (.A1(_22158_),
    .A2(_22161_),
    .A3(_22164_),
    .ZN(_04616_));
 AND3_X1 _27999_ (.A1(_22167_),
    .A2(_04615_),
    .A3(_04616_),
    .ZN(_04617_));
 INV_X1 _28000_ (.A(_22157_),
    .ZN(_04618_));
 NAND3_X1 _28001_ (.A1(_22158_),
    .A2(_22161_),
    .A3(_22164_),
    .ZN(_04619_));
 INV_X1 _28002_ (.A(_22166_),
    .ZN(_04620_));
 AOI21_X1 _28003_ (.A(_22160_),
    .B1(_22163_),
    .B2(_22161_),
    .ZN(_04621_));
 INV_X1 _28004_ (.A(_22158_),
    .ZN(_04622_));
 OAI221_X1 _28005_ (.A(_04618_),
    .B1(_04619_),
    .B2(_04620_),
    .C1(_04621_),
    .C2(_04622_),
    .ZN(_04623_));
 AOI221_X4 _28006_ (.A(_04611_),
    .B1(_04614_),
    .B2(_04617_),
    .C1(_04615_),
    .C2(_04623_),
    .ZN(_04624_));
 AND2_X1 _28007_ (.A1(_22170_),
    .A2(_22173_),
    .ZN(_04625_));
 NAND4_X2 _28008_ (.A1(_22167_),
    .A2(_04615_),
    .A3(_04616_),
    .A4(_04625_),
    .ZN(_04626_));
 NAND2_X2 _28009_ (.A1(_04607_),
    .A2(_04626_),
    .ZN(_04627_));
 OAI22_X1 _28010_ (.A1(_04603_),
    .A2(_04607_),
    .B1(_04624_),
    .B2(_04627_),
    .ZN(_04628_));
 BUF_X4 _28011_ (.A(_04628_),
    .Z(_04629_));
 CLKBUF_X3 _28012_ (.A(_04629_),
    .Z(_04630_));
 OAI21_X1 _28013_ (.A(_04585_),
    .B1(_04589_),
    .B2(_04630_),
    .ZN(_04631_));
 MUX2_X1 _28014_ (.A(\g_reduce0[4].adder.x[15] ),
    .B(\g_reduce0[6].adder.x[15] ),
    .S(_04631_),
    .Z(_00150_));
 INV_X1 _28015_ (.A(_00576_),
    .ZN(_04632_));
 NOR2_X1 _28016_ (.A1(_04632_),
    .A2(_04629_),
    .ZN(_04633_));
 AOI21_X4 _28017_ (.A(_04633_),
    .B1(_04629_),
    .B2(_22174_),
    .ZN(_22266_));
 INV_X1 _28018_ (.A(_22266_),
    .ZN(_22260_));
 MUX2_X2 _28019_ (.A(_22141_),
    .B(_00579_),
    .S(_04629_),
    .Z(_14173_));
 NAND2_X1 _28020_ (.A1(_04593_),
    .A2(_04591_),
    .ZN(_04634_));
 OR2_X1 _28021_ (.A1(_04582_),
    .A2(_22138_),
    .ZN(_04635_));
 OR2_X1 _28022_ (.A1(\g_reduce0[6].adder.x[12] ),
    .A2(_00584_),
    .ZN(_04636_));
 MUX2_X1 _28023_ (.A(_04635_),
    .B(_04636_),
    .S(_04628_),
    .Z(_04637_));
 OR4_X2 _28024_ (.A1(\g_reduce0[6].adder.x[11] ),
    .A2(_00579_),
    .A3(_04624_),
    .A4(_04627_),
    .ZN(_04638_));
 NAND2_X1 _28025_ (.A1(_22178_),
    .A2(_04600_),
    .ZN(_04639_));
 INV_X1 _28026_ (.A(_22175_),
    .ZN(_04640_));
 AOI21_X1 _28027_ (.A(_22142_),
    .B1(_04640_),
    .B2(_04597_),
    .ZN(_04641_));
 OAI221_X2 _28028_ (.A(_04590_),
    .B1(_04606_),
    .B2(_04641_),
    .C1(_04592_),
    .C2(_04594_),
    .ZN(_04642_));
 NAND3_X1 _28029_ (.A1(_04604_),
    .A2(_04597_),
    .A3(_04602_),
    .ZN(_04643_));
 NOR2_X1 _28030_ (.A1(\g_reduce0[6].adder.x[11] ),
    .A2(_00579_),
    .ZN(_04644_));
 NAND4_X2 _28031_ (.A1(_04600_),
    .A2(_04642_),
    .A3(_04643_),
    .A4(_04644_),
    .ZN(_04645_));
 NOR2_X1 _28032_ (.A1(_04581_),
    .A2(_22141_),
    .ZN(_04646_));
 AND2_X1 _28033_ (.A1(_04600_),
    .A2(_04646_),
    .ZN(_04647_));
 OAI221_X2 _28034_ (.A(_04647_),
    .B1(_04627_),
    .B2(_04624_),
    .C1(_04603_),
    .C2(_04607_),
    .ZN(_04648_));
 AND4_X1 _28035_ (.A1(_04638_),
    .A2(_04639_),
    .A3(_04645_),
    .A4(_04648_),
    .ZN(_04649_));
 AOI21_X2 _28036_ (.A(_04634_),
    .B1(_04637_),
    .B2(_04649_),
    .ZN(_04650_));
 NOR2_X1 _28037_ (.A1(\g_reduce0[4].adder.x[13] ),
    .A2(_22135_),
    .ZN(_04651_));
 NOR2_X1 _28038_ (.A1(\g_reduce0[6].adder.x[13] ),
    .A2(_00587_),
    .ZN(_04652_));
 MUX2_X2 _28039_ (.A(_04651_),
    .B(_04652_),
    .S(_04628_),
    .Z(_04653_));
 NOR2_X1 _28040_ (.A1(_04582_),
    .A2(_22138_),
    .ZN(_04654_));
 NOR2_X1 _28041_ (.A1(\g_reduce0[6].adder.x[12] ),
    .A2(_00584_),
    .ZN(_04655_));
 MUX2_X2 _28042_ (.A(_04654_),
    .B(_04655_),
    .S(_04628_),
    .Z(_04656_));
 NAND4_X4 _28043_ (.A1(_04638_),
    .A2(_04639_),
    .A3(_04645_),
    .A4(_04648_),
    .ZN(_04657_));
 NOR4_X4 _28044_ (.A1(_04593_),
    .A2(_04653_),
    .A3(_04656_),
    .A4(_04657_),
    .ZN(_04658_));
 NOR2_X1 _28045_ (.A1(_04593_),
    .A2(_04591_),
    .ZN(_04659_));
 MUX2_X1 _28046_ (.A(_04659_),
    .B(_04593_),
    .S(_04653_),
    .Z(_04660_));
 NOR3_X4 _28047_ (.A1(_04650_),
    .A2(_04658_),
    .A3(_04660_),
    .ZN(_04661_));
 CLKBUF_X3 _28048_ (.A(_04661_),
    .Z(_04662_));
 MUX2_X2 _28049_ (.A(_04646_),
    .B(_04644_),
    .S(_04628_),
    .Z(_04663_));
 NOR3_X4 _28050_ (.A1(_22178_),
    .A2(_04600_),
    .A3(_04663_),
    .ZN(_04664_));
 NOR2_X4 _28051_ (.A1(_04657_),
    .A2(_04664_),
    .ZN(_04665_));
 BUF_X4 _28052_ (.A(_04605_),
    .Z(_04666_));
 BUF_X4 _28053_ (.A(_22179_),
    .Z(_04667_));
 MUX2_X1 _28054_ (.A(_00585_),
    .B(_22144_),
    .S(_04628_),
    .Z(_04668_));
 OAI21_X1 _28055_ (.A(_04666_),
    .B1(_04667_),
    .B2(_04668_),
    .ZN(_04669_));
 MUX2_X1 _28056_ (.A(_00586_),
    .B(_22147_),
    .S(_04628_),
    .Z(_04670_));
 NOR2_X4 _28057_ (.A1(_04666_),
    .A2(_04667_),
    .ZN(_04671_));
 NAND2_X1 _28058_ (.A1(_04670_),
    .A2(_04671_),
    .ZN(_04672_));
 NAND2_X1 _28059_ (.A1(_04669_),
    .A2(_04672_),
    .ZN(_04673_));
 OR2_X1 _28060_ (.A1(_04665_),
    .A2(_04673_),
    .ZN(_04674_));
 MUX2_X1 _28061_ (.A(_00578_),
    .B(_22165_),
    .S(_04628_),
    .Z(_04675_));
 MUX2_X1 _28062_ (.A(_22171_),
    .B(_00575_),
    .S(_04630_),
    .Z(_04676_));
 INV_X2 _28063_ (.A(_04667_),
    .ZN(_04677_));
 MUX2_X1 _28064_ (.A(_04675_),
    .B(_04676_),
    .S(_04677_),
    .Z(_04678_));
 MUX2_X1 _28065_ (.A(_00577_),
    .B(_22162_),
    .S(_04630_),
    .Z(_04679_));
 MUX2_X1 _28066_ (.A(_00574_),
    .B(_22168_),
    .S(_04630_),
    .Z(_04680_));
 MUX2_X1 _28067_ (.A(_04679_),
    .B(_04680_),
    .S(_04677_),
    .Z(_04681_));
 MUX2_X1 _28068_ (.A(_04678_),
    .B(_04681_),
    .S(_04666_),
    .Z(_04682_));
 MUX2_X1 _28069_ (.A(_00583_),
    .B(_22153_),
    .S(_04630_),
    .Z(_04683_));
 MUX2_X1 _28070_ (.A(_00582_),
    .B(_22150_),
    .S(_04630_),
    .Z(_04684_));
 MUX2_X1 _28071_ (.A(_04683_),
    .B(_04684_),
    .S(_04666_),
    .Z(_04685_));
 MUX2_X1 _28072_ (.A(_00581_),
    .B(_22159_),
    .S(_04630_),
    .Z(_04686_));
 MUX2_X1 _28073_ (.A(_00580_),
    .B(_22156_),
    .S(_04630_),
    .Z(_04687_));
 MUX2_X1 _28074_ (.A(_04686_),
    .B(_04687_),
    .S(_04666_),
    .Z(_04688_));
 MUX2_X1 _28075_ (.A(_04685_),
    .B(_04688_),
    .S(_04677_),
    .Z(_04689_));
 MUX2_X1 _28076_ (.A(_04682_),
    .B(_04689_),
    .S(_04665_),
    .Z(_04690_));
 NAND4_X1 _28077_ (.A1(_04632_),
    .A2(_22174_),
    .A3(_04642_),
    .A4(_04643_),
    .ZN(_04691_));
 NAND4_X1 _28078_ (.A1(_04632_),
    .A2(_22174_),
    .A3(_04607_),
    .A4(_04626_),
    .ZN(_04692_));
 OR2_X1 _28079_ (.A1(_04624_),
    .A2(_04692_),
    .ZN(_04693_));
 NOR2_X1 _28080_ (.A1(_04632_),
    .A2(_22174_),
    .ZN(_04694_));
 OAI221_X1 _28081_ (.A(_04694_),
    .B1(_04627_),
    .B2(_04624_),
    .C1(_04603_),
    .C2(_04607_),
    .ZN(_04695_));
 AND3_X2 _28082_ (.A1(_04691_),
    .A2(_04693_),
    .A3(_04695_),
    .ZN(_22177_));
 OR4_X2 _28083_ (.A1(_04591_),
    .A2(_04656_),
    .A3(_04663_),
    .A4(_22177_),
    .ZN(_04696_));
 AND2_X1 _28084_ (.A1(_04597_),
    .A2(_04601_),
    .ZN(_04697_));
 AOI22_X4 _28085_ (.A1(_04601_),
    .A2(_04663_),
    .B1(_22177_),
    .B2(_04697_),
    .ZN(_04698_));
 OR4_X2 _28086_ (.A1(_04591_),
    .A2(_04597_),
    .A3(_04656_),
    .A4(_04663_),
    .ZN(_04699_));
 INV_X1 _28087_ (.A(_04591_),
    .ZN(_04700_));
 OR2_X1 _28088_ (.A1(_04591_),
    .A2(_04600_),
    .ZN(_04701_));
 MUX2_X2 _28089_ (.A(_04700_),
    .B(_04701_),
    .S(_04637_),
    .Z(_04702_));
 NAND4_X4 _28090_ (.A1(_04696_),
    .A2(_04698_),
    .A3(_04699_),
    .A4(_04702_),
    .ZN(_04703_));
 MUX2_X1 _28091_ (.A(_04674_),
    .B(_04690_),
    .S(_04703_),
    .Z(_04704_));
 OR2_X1 _28092_ (.A1(_04662_),
    .A2(_04704_),
    .ZN(_22246_));
 INV_X1 _28093_ (.A(_22246_),
    .ZN(_22243_));
 AOI21_X1 _28094_ (.A(_04667_),
    .B1(_04668_),
    .B2(_04604_),
    .ZN(_04705_));
 INV_X1 _28095_ (.A(_04705_),
    .ZN(_04706_));
 MUX2_X1 _28096_ (.A(_04686_),
    .B(_04675_),
    .S(_04677_),
    .Z(_04707_));
 MUX2_X1 _28097_ (.A(_04681_),
    .B(_04707_),
    .S(_04666_),
    .Z(_04708_));
 MUX2_X1 _28098_ (.A(_04706_),
    .B(_04708_),
    .S(_04703_),
    .Z(_04709_));
 MUX2_X1 _28099_ (.A(_04670_),
    .B(_04683_),
    .S(_04677_),
    .Z(_04710_));
 MUX2_X1 _28100_ (.A(_04684_),
    .B(_04687_),
    .S(_04677_),
    .Z(_04711_));
 MUX2_X1 _28101_ (.A(_04710_),
    .B(_04711_),
    .S(_04604_),
    .Z(_04712_));
 NAND2_X1 _28102_ (.A1(_04665_),
    .A2(_04703_),
    .ZN(_04713_));
 OAI22_X1 _28103_ (.A1(_04665_),
    .A2(_04709_),
    .B1(_04712_),
    .B2(_04713_),
    .ZN(_04714_));
 INV_X1 _28104_ (.A(_04714_),
    .ZN(_04715_));
 OR2_X1 _28105_ (.A1(_04662_),
    .A2(_04715_),
    .ZN(_14169_));
 INV_X1 _28106_ (.A(_14169_),
    .ZN(_14164_));
 AND4_X1 _28107_ (.A1(_04696_),
    .A2(_04698_),
    .A3(_04699_),
    .A4(_04702_),
    .ZN(_04716_));
 BUF_X4 _28108_ (.A(_04716_),
    .Z(_04717_));
 OR2_X1 _28109_ (.A1(_04662_),
    .A2(_04717_),
    .ZN(_04718_));
 BUF_X2 _28110_ (.A(_04718_),
    .Z(_04719_));
 NOR2_X1 _28111_ (.A1(_04665_),
    .A2(_04719_),
    .ZN(_04720_));
 NAND2_X1 _28112_ (.A1(_04705_),
    .A2(_04720_),
    .ZN(_22198_));
 INV_X1 _28113_ (.A(_22198_),
    .ZN(_22202_));
 OR2_X1 _28114_ (.A1(_04674_),
    .A2(_04719_),
    .ZN(_22192_));
 INV_X1 _28115_ (.A(_22192_),
    .ZN(_22195_));
 AND2_X1 _28116_ (.A1(_00582_),
    .A2(_04671_),
    .ZN(_04721_));
 AND2_X1 _28117_ (.A1(_22150_),
    .A2(_04671_),
    .ZN(_04722_));
 MUX2_X1 _28118_ (.A(_04721_),
    .B(_04722_),
    .S(_04628_),
    .Z(_04723_));
 NAND2_X2 _28119_ (.A1(_04604_),
    .A2(_04667_),
    .ZN(_04724_));
 INV_X1 _28120_ (.A(_04724_),
    .ZN(_04725_));
 NOR2_X2 _28121_ (.A1(_04604_),
    .A2(_04667_),
    .ZN(_04726_));
 AOI221_X2 _28122_ (.A(_04723_),
    .B1(_04725_),
    .B2(_04668_),
    .C1(_04670_),
    .C2(_04726_),
    .ZN(_04727_));
 NAND2_X1 _28123_ (.A1(_04720_),
    .A2(_04727_),
    .ZN(_22226_));
 INV_X1 _28124_ (.A(_22226_),
    .ZN(_22230_));
 MUX2_X1 _28125_ (.A(_04670_),
    .B(_04668_),
    .S(_04666_),
    .Z(_04728_));
 MUX2_X1 _28126_ (.A(_04685_),
    .B(_04728_),
    .S(_04667_),
    .Z(_04729_));
 NAND2_X1 _28127_ (.A1(_04604_),
    .A2(_04677_),
    .ZN(_04730_));
 MUX2_X1 _28128_ (.A(_04729_),
    .B(_04730_),
    .S(_04665_),
    .Z(_04731_));
 OR2_X1 _28129_ (.A1(_04719_),
    .A2(_04731_),
    .ZN(_22206_));
 INV_X1 _28130_ (.A(_22206_),
    .ZN(_22209_));
 MUX2_X1 _28131_ (.A(_04712_),
    .B(_04706_),
    .S(_04665_),
    .Z(_04732_));
 NOR2_X1 _28132_ (.A1(_04719_),
    .A2(_04732_),
    .ZN(_22213_));
 INV_X1 _28133_ (.A(_22213_),
    .ZN(_22216_));
 MUX2_X1 _28134_ (.A(_04689_),
    .B(_04673_),
    .S(_04665_),
    .Z(_04733_));
 NOR2_X1 _28135_ (.A1(_04719_),
    .A2(_04733_),
    .ZN(_22219_));
 INV_X1 _28136_ (.A(_22219_),
    .ZN(_22223_));
 NAND2_X2 _28137_ (.A1(_04666_),
    .A2(_04677_),
    .ZN(_04734_));
 OAI22_X1 _28138_ (.A1(_00580_),
    .A2(_04724_),
    .B1(_04734_),
    .B2(_00581_),
    .ZN(_04735_));
 NAND2_X1 _28139_ (.A1(_04666_),
    .A2(_04667_),
    .ZN(_04736_));
 OAI22_X1 _28140_ (.A1(_00577_),
    .A2(_04730_),
    .B1(_04736_),
    .B2(_00583_),
    .ZN(_04737_));
 NOR2_X1 _28141_ (.A1(_04735_),
    .A2(_04737_),
    .ZN(_04738_));
 OAI22_X1 _28142_ (.A1(_22156_),
    .A2(_04724_),
    .B1(_04734_),
    .B2(_22159_),
    .ZN(_04739_));
 OAI22_X1 _28143_ (.A1(_22162_),
    .A2(_04730_),
    .B1(_04736_),
    .B2(_22153_),
    .ZN(_04740_));
 NOR2_X1 _28144_ (.A1(_04739_),
    .A2(_04740_),
    .ZN(_04741_));
 MUX2_X1 _28145_ (.A(_04738_),
    .B(_04741_),
    .S(_04629_),
    .Z(_04742_));
 AOI21_X1 _28146_ (.A(_04721_),
    .B1(_04726_),
    .B2(_00586_),
    .ZN(_04743_));
 AOI21_X1 _28147_ (.A(_04722_),
    .B1(_04726_),
    .B2(_22147_),
    .ZN(_04744_));
 MUX2_X1 _28148_ (.A(_04743_),
    .B(_04744_),
    .S(_04629_),
    .Z(_04745_));
 INV_X1 _28149_ (.A(_00585_),
    .ZN(_04746_));
 INV_X1 _28150_ (.A(_22144_),
    .ZN(_04747_));
 MUX2_X1 _28151_ (.A(_04746_),
    .B(_04747_),
    .S(_04629_),
    .Z(_04748_));
 OAI21_X1 _28152_ (.A(_04745_),
    .B1(_04724_),
    .B2(_04748_),
    .ZN(_04749_));
 MUX2_X1 _28153_ (.A(_04742_),
    .B(_04749_),
    .S(_04665_),
    .Z(_04750_));
 NOR2_X1 _28154_ (.A1(_04719_),
    .A2(_04750_),
    .ZN(_22237_));
 INV_X1 _28155_ (.A(_22237_),
    .ZN(_22240_));
 MUX2_X1 _28156_ (.A(_04687_),
    .B(_04679_),
    .S(_04677_),
    .Z(_04751_));
 MUX2_X1 _28157_ (.A(_04707_),
    .B(_04751_),
    .S(_04666_),
    .Z(_04752_));
 MUX2_X1 _28158_ (.A(_04730_),
    .B(_04752_),
    .S(_04703_),
    .Z(_04753_));
 NOR2_X1 _28159_ (.A1(_04665_),
    .A2(_04753_),
    .ZN(_04754_));
 NOR2_X1 _28160_ (.A1(_04713_),
    .A2(_04729_),
    .ZN(_04755_));
 NOR2_X1 _28161_ (.A1(_04754_),
    .A2(_04755_),
    .ZN(_04756_));
 OR2_X1 _28162_ (.A1(_04662_),
    .A2(_04756_),
    .ZN(_22233_));
 INV_X1 _28163_ (.A(_22233_),
    .ZN(_22187_));
 INV_X1 _28164_ (.A(_22200_),
    .ZN(_04757_));
 INV_X1 _28165_ (.A(_22193_),
    .ZN(_04758_));
 NAND2_X1 _28166_ (.A1(_04757_),
    .A2(_04758_),
    .ZN(_04759_));
 INV_X1 _28167_ (.A(_22228_),
    .ZN(_04760_));
 OR3_X1 _28168_ (.A1(_22217_),
    .A2(_22207_),
    .A3(_22224_),
    .ZN(_04761_));
 INV_X1 _28169_ (.A(_22241_),
    .ZN(_04762_));
 AOI21_X1 _28170_ (.A(_22234_),
    .B1(_14171_),
    .B2(_22235_),
    .ZN(_04763_));
 CLKBUF_X2 _28171_ (.A(_22239_),
    .Z(_04764_));
 OAI21_X1 _28172_ (.A(_04762_),
    .B1(_04763_),
    .B2(_04764_),
    .ZN(_04765_));
 BUF_X2 _28173_ (.A(_22222_),
    .Z(_04766_));
 INV_X1 _28174_ (.A(_04766_),
    .ZN(_04767_));
 AOI21_X1 _28175_ (.A(_04761_),
    .B1(_04765_),
    .B2(_04767_),
    .ZN(_04768_));
 BUF_X2 _28176_ (.A(_22229_),
    .Z(_04769_));
 INV_X1 _28177_ (.A(_22208_),
    .ZN(_04770_));
 INV_X1 _28178_ (.A(_22217_),
    .ZN(_04771_));
 AOI21_X1 _28179_ (.A(_04770_),
    .B1(_04771_),
    .B2(_22215_),
    .ZN(_04772_));
 OAI21_X1 _28180_ (.A(_04769_),
    .B1(_22207_),
    .B2(_04772_),
    .ZN(_04773_));
 OAI21_X1 _28181_ (.A(_04760_),
    .B1(_04768_),
    .B2(_04773_),
    .ZN(_04774_));
 BUF_X2 _28182_ (.A(_22194_),
    .Z(_04775_));
 AOI21_X1 _28183_ (.A(_04759_),
    .B1(_04774_),
    .B2(_04775_),
    .ZN(_04776_));
 INV_X1 _28184_ (.A(\g_reduce0[6].adder.x[15] ),
    .ZN(_04777_));
 NOR2_X2 _28185_ (.A1(_04777_),
    .A2(\g_reduce0[4].adder.x[15] ),
    .ZN(_04778_));
 AND2_X1 _28186_ (.A1(_04777_),
    .A2(\g_reduce0[4].adder.x[15] ),
    .ZN(_04779_));
 OR2_X1 _28187_ (.A1(_04778_),
    .A2(_04779_),
    .ZN(_04780_));
 BUF_X4 _28188_ (.A(_04780_),
    .Z(_04781_));
 MUX2_X2 _28189_ (.A(_22203_),
    .B(_04776_),
    .S(_04781_),
    .Z(_04782_));
 INV_X2 _28190_ (.A(_22201_),
    .ZN(_04783_));
 XNOR2_X2 _28191_ (.A(\g_reduce0[6].adder.x[15] ),
    .B(\g_reduce0[4].adder.x[15] ),
    .ZN(_04784_));
 BUF_X4 _28192_ (.A(_04784_),
    .Z(_04785_));
 OAI21_X2 _28193_ (.A(_04783_),
    .B1(_04757_),
    .B2(_04785_),
    .ZN(_04786_));
 INV_X1 _28194_ (.A(_22231_),
    .ZN(_04787_));
 OR2_X1 _28195_ (.A1(_22210_),
    .A2(_22214_),
    .ZN(_04788_));
 NOR2_X1 _28196_ (.A1(_22221_),
    .A2(_22238_),
    .ZN(_04789_));
 BUF_X1 _28197_ (.A(_22190_),
    .Z(_04790_));
 AOI21_X2 _28198_ (.A(_22189_),
    .B1(_14167_),
    .B2(_04790_),
    .ZN(_04791_));
 INV_X2 _28199_ (.A(_04764_),
    .ZN(_04792_));
 OAI21_X1 _28200_ (.A(_04789_),
    .B1(_04791_),
    .B2(_04792_),
    .ZN(_04793_));
 INV_X1 _28201_ (.A(_22215_),
    .ZN(_04794_));
 INV_X1 _28202_ (.A(_22221_),
    .ZN(_04795_));
 AOI21_X2 _28203_ (.A(_04794_),
    .B1(_04767_),
    .B2(_04795_),
    .ZN(_04796_));
 AOI21_X1 _28204_ (.A(_04788_),
    .B1(_04793_),
    .B2(_04796_),
    .ZN(_04797_));
 INV_X1 _28205_ (.A(_04769_),
    .ZN(_04798_));
 OAI21_X1 _28206_ (.A(_04798_),
    .B1(_22210_),
    .B2(_04770_),
    .ZN(_04799_));
 OAI21_X1 _28207_ (.A(_04787_),
    .B1(_04797_),
    .B2(_04799_),
    .ZN(_04800_));
 INV_X1 _28208_ (.A(_04775_),
    .ZN(_04801_));
 AOI21_X2 _28209_ (.A(_22196_),
    .B1(_04800_),
    .B2(_04801_),
    .ZN(_04802_));
 AOI21_X4 _28210_ (.A(_04786_),
    .B1(_04802_),
    .B2(_04785_),
    .ZN(_04803_));
 NOR2_X4 _28211_ (.A1(_04782_),
    .A2(_04803_),
    .ZN(_04804_));
 INV_X1 _28212_ (.A(_22224_),
    .ZN(_04805_));
 NAND3_X1 _28213_ (.A1(_04771_),
    .A2(_04805_),
    .A3(_04762_),
    .ZN(_04806_));
 INV_X1 _28214_ (.A(_22234_),
    .ZN(_04807_));
 INV_X1 _28215_ (.A(_22235_),
    .ZN(_04808_));
 AOI21_X1 _28216_ (.A(_22185_),
    .B1(_14170_),
    .B2(_22186_),
    .ZN(_04809_));
 OAI21_X2 _28217_ (.A(_04807_),
    .B1(_04808_),
    .B2(_04809_),
    .ZN(_04810_));
 AOI21_X2 _28218_ (.A(_04806_),
    .B1(_04810_),
    .B2(_04792_),
    .ZN(_04811_));
 AOI21_X1 _28219_ (.A(_22215_),
    .B1(_04766_),
    .B2(_04805_),
    .ZN(_04812_));
 OAI21_X1 _28220_ (.A(_22208_),
    .B1(_22217_),
    .B2(_04812_),
    .ZN(_04813_));
 NAND2_X1 _28221_ (.A1(_04775_),
    .A2(_04769_),
    .ZN(_04814_));
 OR3_X1 _28222_ (.A1(_04811_),
    .A2(_04813_),
    .A3(_04814_),
    .ZN(_04815_));
 AOI21_X1 _28223_ (.A(_22228_),
    .B1(_22207_),
    .B2(_04769_),
    .ZN(_04816_));
 INV_X1 _28224_ (.A(_04816_),
    .ZN(_04817_));
 AOI21_X1 _28225_ (.A(_22193_),
    .B1(_04817_),
    .B2(_04775_),
    .ZN(_04818_));
 AOI21_X2 _28226_ (.A(_04783_),
    .B1(_04815_),
    .B2(_04818_),
    .ZN(_04819_));
 OAI21_X4 _28227_ (.A(_04781_),
    .B1(_04819_),
    .B2(_22200_),
    .ZN(_04820_));
 NOR2_X1 _28228_ (.A1(_04804_),
    .A2(_04820_),
    .ZN(_04821_));
 AOI21_X1 _28229_ (.A(_04775_),
    .B1(_04769_),
    .B2(_04787_),
    .ZN(_04822_));
 NOR2_X1 _28230_ (.A1(_22196_),
    .A2(_04822_),
    .ZN(_04823_));
 NOR3_X1 _28231_ (.A1(_22231_),
    .A2(_22196_),
    .A3(_22210_),
    .ZN(_04824_));
 INV_X1 _28232_ (.A(_22189_),
    .ZN(_04825_));
 AOI21_X2 _28233_ (.A(_22183_),
    .B1(_14166_),
    .B2(_22184_),
    .ZN(_04826_));
 NAND2_X1 _28234_ (.A1(_04764_),
    .A2(_04790_),
    .ZN(_04827_));
 OAI22_X2 _28235_ (.A1(_04825_),
    .A2(_04792_),
    .B1(_04826_),
    .B2(_04827_),
    .ZN(_04828_));
 OR3_X1 _28236_ (.A1(_22214_),
    .A2(_22221_),
    .A3(_22238_),
    .ZN(_04829_));
 OAI221_X2 _28237_ (.A(_04770_),
    .B1(_22214_),
    .B2(_04796_),
    .C1(_04828_),
    .C2(_04829_),
    .ZN(_04830_));
 AOI21_X2 _28238_ (.A(_04823_),
    .B1(_04824_),
    .B2(_04830_),
    .ZN(_04831_));
 AOI21_X2 _28239_ (.A(_22203_),
    .B1(_04783_),
    .B2(_04831_),
    .ZN(_04832_));
 NOR2_X2 _28240_ (.A1(_04781_),
    .A2(_04832_),
    .ZN(_04833_));
 OR2_X2 _28241_ (.A1(_04782_),
    .A2(_04803_),
    .ZN(_04834_));
 NOR2_X1 _28242_ (.A1(_04833_),
    .A2(_04834_),
    .ZN(_04835_));
 OAI21_X4 _28243_ (.A(_04671_),
    .B1(_04664_),
    .B2(_04657_),
    .ZN(_04836_));
 OR3_X4 _28244_ (.A1(_04661_),
    .A2(_04717_),
    .A3(_04836_),
    .ZN(_04837_));
 MUX2_X2 _28245_ (.A(_04821_),
    .B(_04835_),
    .S(_04837_),
    .Z(_04838_));
 NAND2_X1 _28246_ (.A1(_04781_),
    .A2(_04774_),
    .ZN(_04839_));
 OR2_X1 _28247_ (.A1(_04781_),
    .A2(_04800_),
    .ZN(_04840_));
 AND3_X2 _28248_ (.A1(_04775_),
    .A2(_04839_),
    .A3(_04840_),
    .ZN(_04841_));
 AOI21_X4 _28249_ (.A(_04775_),
    .B1(_04839_),
    .B2(_04840_),
    .ZN(_04842_));
 NAND2_X1 _28250_ (.A1(_22210_),
    .A2(_04785_),
    .ZN(_04843_));
 MUX2_X1 _28251_ (.A(_22207_),
    .B(_04830_),
    .S(_04784_),
    .Z(_04844_));
 NOR2_X1 _28252_ (.A1(_04811_),
    .A2(_04813_),
    .ZN(_04845_));
 OAI21_X2 _28253_ (.A(_04843_),
    .B1(_04844_),
    .B2(_04845_),
    .ZN(_04846_));
 XNOR2_X2 _28254_ (.A(_04798_),
    .B(_04846_),
    .ZN(_04847_));
 AOI21_X1 _28255_ (.A(_22214_),
    .B1(_04796_),
    .B2(_04793_),
    .ZN(_04848_));
 OR2_X1 _28256_ (.A1(_04780_),
    .A2(_04848_),
    .ZN(_04849_));
 AOI21_X1 _28257_ (.A(_22224_),
    .B1(_04765_),
    .B2(_04767_),
    .ZN(_04850_));
 OAI221_X2 _28258_ (.A(_04771_),
    .B1(_04778_),
    .B2(_04779_),
    .C1(_04850_),
    .C2(_22215_),
    .ZN(_04851_));
 AOI21_X1 _28259_ (.A(_04770_),
    .B1(_04849_),
    .B2(_04851_),
    .ZN(_04852_));
 AND3_X1 _28260_ (.A1(_04770_),
    .A2(_04849_),
    .A3(_04851_),
    .ZN(_04853_));
 INV_X1 _28261_ (.A(_22238_),
    .ZN(_04854_));
 OAI221_X1 _28262_ (.A(_04854_),
    .B1(_04826_),
    .B2(_04827_),
    .C1(_04792_),
    .C2(_04825_),
    .ZN(_04855_));
 AOI21_X1 _28263_ (.A(_22221_),
    .B1(_04855_),
    .B2(_04766_),
    .ZN(_04856_));
 OR2_X1 _28264_ (.A1(_04780_),
    .A2(_04856_),
    .ZN(_04857_));
 AOI21_X1 _28265_ (.A(_22241_),
    .B1(_04810_),
    .B2(_04792_),
    .ZN(_04858_));
 OAI221_X2 _28266_ (.A(_04805_),
    .B1(_04778_),
    .B2(_04779_),
    .C1(_04858_),
    .C2(_04766_),
    .ZN(_04859_));
 AND3_X1 _28267_ (.A1(_04794_),
    .A2(_04857_),
    .A3(_04859_),
    .ZN(_04860_));
 AOI21_X2 _28268_ (.A(_04794_),
    .B1(_04857_),
    .B2(_04859_),
    .ZN(_04861_));
 OR4_X1 _28269_ (.A1(_04852_),
    .A2(_04853_),
    .A3(_04860_),
    .A4(_04861_),
    .ZN(_04862_));
 AOI211_X2 _28270_ (.A(_04841_),
    .B(_04842_),
    .C1(_04847_),
    .C2(_04862_),
    .ZN(_04863_));
 NOR3_X1 _28271_ (.A1(_04811_),
    .A2(_04813_),
    .A3(_04814_),
    .ZN(_04864_));
 OAI21_X1 _28272_ (.A(_04758_),
    .B1(_04816_),
    .B2(_04801_),
    .ZN(_04865_));
 NOR2_X1 _28273_ (.A1(_04864_),
    .A2(_04865_),
    .ZN(_04866_));
 MUX2_X2 _28274_ (.A(_04831_),
    .B(_04866_),
    .S(_04781_),
    .Z(_04867_));
 XNOR2_X2 _28275_ (.A(_22201_),
    .B(_04867_),
    .ZN(_04868_));
 OR2_X2 _28276_ (.A1(_04863_),
    .A2(_04868_),
    .ZN(_04869_));
 OAI211_X2 _28277_ (.A(_04671_),
    .B(_04820_),
    .C1(_04657_),
    .C2(_04664_),
    .ZN(_04870_));
 OAI33_X1 _28278_ (.A1(_04778_),
    .A2(_04779_),
    .A3(_04832_),
    .B1(_04870_),
    .B2(_04662_),
    .B3(_04717_),
    .ZN(_04871_));
 BUF_X4 _28279_ (.A(_04871_),
    .Z(_04872_));
 NOR2_X4 _28280_ (.A1(_04869_),
    .A2(_04872_),
    .ZN(_04873_));
 OR2_X1 _28281_ (.A1(_04852_),
    .A2(_04853_),
    .ZN(_04874_));
 BUF_X1 _28282_ (.A(_04874_),
    .Z(_04875_));
 NOR2_X1 _28283_ (.A1(_04784_),
    .A2(_04765_),
    .ZN(_04876_));
 OAI21_X2 _28284_ (.A(_04854_),
    .B1(_04791_),
    .B2(_04792_),
    .ZN(_04877_));
 AOI21_X4 _28285_ (.A(_04876_),
    .B1(_04877_),
    .B2(_04785_),
    .ZN(_04878_));
 XNOR2_X2 _28286_ (.A(_04766_),
    .B(_04878_),
    .ZN(_04879_));
 NOR4_X1 _28287_ (.A1(_04841_),
    .A2(_04842_),
    .A3(_04875_),
    .A4(_04879_),
    .ZN(_04880_));
 INV_X1 _28288_ (.A(_04790_),
    .ZN(_04881_));
 OAI21_X1 _28289_ (.A(_04825_),
    .B1(_04881_),
    .B2(_04826_),
    .ZN(_04882_));
 NAND2_X1 _28290_ (.A1(_04784_),
    .A2(_04882_),
    .ZN(_04883_));
 OAI21_X2 _28291_ (.A(_04883_),
    .B1(_04810_),
    .B2(_04784_),
    .ZN(_04884_));
 XNOR2_X2 _28292_ (.A(_04764_),
    .B(_04884_),
    .ZN(_04885_));
 MUX2_X2 _28293_ (.A(_14172_),
    .B(_14168_),
    .S(_04785_),
    .Z(_04886_));
 XOR2_X1 _28294_ (.A(_14171_),
    .B(_22235_),
    .Z(_04887_));
 XOR2_X1 _28295_ (.A(_14167_),
    .B(_04790_),
    .Z(_04888_));
 MUX2_X1 _28296_ (.A(_04887_),
    .B(_04888_),
    .S(_04784_),
    .Z(_04889_));
 CLKBUF_X3 _28297_ (.A(_04889_),
    .Z(_04890_));
 OAI21_X2 _28298_ (.A(_04885_),
    .B1(_04886_),
    .B2(_04890_),
    .ZN(_04891_));
 INV_X1 _28299_ (.A(_04891_),
    .ZN(_04892_));
 MUX2_X2 _28300_ (.A(_22247_),
    .B(_22245_),
    .S(_04784_),
    .Z(_04893_));
 NOR2_X1 _28301_ (.A1(_04890_),
    .A2(_04893_),
    .ZN(_04894_));
 NAND2_X2 _28302_ (.A1(_04785_),
    .A2(_04894_),
    .ZN(_04895_));
 OR2_X2 _28303_ (.A1(_04662_),
    .A2(_04895_),
    .ZN(_04896_));
 OAI21_X2 _28304_ (.A(_04727_),
    .B1(_04664_),
    .B2(_04657_),
    .ZN(_04897_));
 NOR2_X1 _28305_ (.A1(_04675_),
    .A2(_04736_),
    .ZN(_04898_));
 OAI221_X2 _28306_ (.A(_04629_),
    .B1(_04724_),
    .B2(_22168_),
    .C1(_04734_),
    .C2(_00575_),
    .ZN(_04899_));
 OAI22_X1 _28307_ (.A1(_00574_),
    .A2(_04724_),
    .B1(_04734_),
    .B2(_22171_),
    .ZN(_04900_));
 OR2_X1 _28308_ (.A1(_04629_),
    .A2(_04900_),
    .ZN(_04901_));
 AND2_X1 _28309_ (.A1(_04899_),
    .A2(_04901_),
    .ZN(_04902_));
 OAI22_X4 _28310_ (.A1(_04657_),
    .A2(_04664_),
    .B1(_04898_),
    .B2(_04902_),
    .ZN(_04903_));
 MUX2_X2 _28311_ (.A(_04897_),
    .B(_04903_),
    .S(_04703_),
    .Z(_04904_));
 OAI21_X2 _28312_ (.A(_04892_),
    .B1(_04896_),
    .B2(_04904_),
    .ZN(_04905_));
 NOR3_X2 _28313_ (.A1(_22247_),
    .A2(_04785_),
    .A3(_04890_),
    .ZN(_04906_));
 OR3_X2 _28314_ (.A1(_04657_),
    .A2(_04664_),
    .A3(_04742_),
    .ZN(_04907_));
 NAND4_X2 _28315_ (.A1(_04703_),
    .A2(_04906_),
    .A3(_04903_),
    .A4(_04907_),
    .ZN(_04908_));
 OR4_X2 _28316_ (.A1(_04661_),
    .A2(_04717_),
    .A3(_04907_),
    .A4(_04895_),
    .ZN(_04909_));
 NAND2_X1 _28317_ (.A1(_04781_),
    .A2(_04894_),
    .ZN(_04910_));
 AOI21_X4 _28318_ (.A(_04662_),
    .B1(_04717_),
    .B2(_04897_),
    .ZN(_04911_));
 OAI211_X4 _28319_ (.A(_04908_),
    .B(_04909_),
    .C1(_04910_),
    .C2(_04911_),
    .ZN(_04912_));
 OAI21_X1 _28320_ (.A(_04880_),
    .B1(_04905_),
    .B2(_04912_),
    .ZN(_04913_));
 AOI21_X1 _28321_ (.A(_04838_),
    .B1(_04873_),
    .B2(_04913_),
    .ZN(_22249_));
 INV_X2 _28322_ (.A(_22249_),
    .ZN(_22251_));
 CLKBUF_X3 _28323_ (.A(_22254_),
    .Z(_04914_));
 INV_X1 _28324_ (.A(_04914_),
    .ZN(_04915_));
 OR2_X2 _28325_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04916_));
 INV_X1 _28326_ (.A(_04890_),
    .ZN(_04917_));
 XNOR2_X2 _28327_ (.A(_04767_),
    .B(_04878_),
    .ZN(_04918_));
 NAND4_X4 _28328_ (.A1(_04916_),
    .A2(_04917_),
    .A3(_04885_),
    .A4(_04918_),
    .ZN(_04919_));
 NOR2_X2 _28329_ (.A1(_04841_),
    .A2(_04842_),
    .ZN(_04920_));
 XNOR2_X2 _28330_ (.A(_04783_),
    .B(_04867_),
    .ZN(_04921_));
 XNOR2_X2 _28331_ (.A(_04769_),
    .B(_04846_),
    .ZN(_04922_));
 NOR2_X1 _28332_ (.A1(_04922_),
    .A2(_04875_),
    .ZN(_04923_));
 AND3_X1 _28333_ (.A1(_04920_),
    .A2(_04921_),
    .A3(_04923_),
    .ZN(_04924_));
 NAND2_X1 _28334_ (.A1(_04919_),
    .A2(_04924_),
    .ZN(_04925_));
 NOR2_X1 _28335_ (.A1(_04834_),
    .A2(_04820_),
    .ZN(_04926_));
 NOR2_X1 _28336_ (.A1(_04833_),
    .A2(_04804_),
    .ZN(_04927_));
 MUX2_X1 _28337_ (.A(_04926_),
    .B(_04927_),
    .S(_04837_),
    .Z(_04928_));
 BUF_X4 _28338_ (.A(_04928_),
    .Z(_04929_));
 AOI21_X4 _28339_ (.A(_04915_),
    .B1(_04925_),
    .B2(_04929_),
    .ZN(_04930_));
 AND4_X1 _28340_ (.A1(_04920_),
    .A2(_04921_),
    .A3(_04919_),
    .A4(_04923_),
    .ZN(_04931_));
 OAI21_X1 _28341_ (.A(_22201_),
    .B1(_04864_),
    .B2(_04865_),
    .ZN(_04932_));
 AOI21_X1 _28342_ (.A(_04785_),
    .B1(_04932_),
    .B2(_04757_),
    .ZN(_04933_));
 NAND2_X1 _28343_ (.A1(_04804_),
    .A2(_04933_),
    .ZN(_04934_));
 OR2_X1 _28344_ (.A1(_04833_),
    .A2(_04804_),
    .ZN(_04935_));
 MUX2_X2 _28345_ (.A(_04934_),
    .B(_04935_),
    .S(_04837_),
    .Z(_04936_));
 NOR3_X4 _28346_ (.A1(_04914_),
    .A2(_04931_),
    .A3(_04936_),
    .ZN(_04937_));
 NOR2_X4 _28347_ (.A1(_04930_),
    .A2(_04937_),
    .ZN(_04938_));
 INV_X4 _28348_ (.A(_04938_),
    .ZN(_22275_));
 XNOR2_X1 _28349_ (.A(_04914_),
    .B(_04931_),
    .ZN(_04939_));
 AND2_X2 _28350_ (.A1(_04929_),
    .A2(_04939_),
    .ZN(_04940_));
 INV_X1 _28351_ (.A(_04919_),
    .ZN(_04941_));
 NOR2_X2 _28352_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04942_));
 XNOR2_X2 _28353_ (.A(_04792_),
    .B(_04884_),
    .ZN(_04943_));
 AND2_X1 _28354_ (.A1(_14168_),
    .A2(_04784_),
    .ZN(_04944_));
 AOI21_X4 _28355_ (.A(_04944_),
    .B1(_04781_),
    .B2(_14172_),
    .ZN(_04945_));
 NOR2_X1 _28356_ (.A1(_04893_),
    .A2(_04945_),
    .ZN(_04946_));
 NOR3_X2 _28357_ (.A1(_04890_),
    .A2(_04943_),
    .A3(_04946_),
    .ZN(_04947_));
 NOR3_X4 _28358_ (.A1(_04942_),
    .A2(_04879_),
    .A3(_04947_),
    .ZN(_04948_));
 CLKBUF_X3 _28359_ (.A(_04863_),
    .Z(_04949_));
 NOR2_X2 _28360_ (.A1(_04949_),
    .A2(_04880_),
    .ZN(_04950_));
 OR4_X1 _28361_ (.A1(_04942_),
    .A2(_04891_),
    .A3(_04879_),
    .A4(_04947_),
    .ZN(_04951_));
 OR2_X1 _28362_ (.A1(_04949_),
    .A2(_04951_),
    .ZN(_04952_));
 NOR2_X1 _28363_ (.A1(_04662_),
    .A2(_04895_),
    .ZN(_04953_));
 OR3_X1 _28364_ (.A1(_22178_),
    .A2(_04600_),
    .A3(_04663_),
    .ZN(_04954_));
 AOI21_X1 _28365_ (.A(_04749_),
    .B1(_04954_),
    .B2(_04649_),
    .ZN(_04955_));
 OR2_X1 _28366_ (.A1(_04675_),
    .A2(_04736_),
    .ZN(_04956_));
 NAND2_X1 _28367_ (.A1(_04899_),
    .A2(_04901_),
    .ZN(_04957_));
 AOI22_X1 _28368_ (.A1(_04649_),
    .A2(_04954_),
    .B1(_04956_),
    .B2(_04957_),
    .ZN(_04958_));
 MUX2_X1 _28369_ (.A(_04955_),
    .B(_04958_),
    .S(_04703_),
    .Z(_04959_));
 AOI21_X1 _28370_ (.A(_04952_),
    .B1(_04953_),
    .B2(_04959_),
    .ZN(_04960_));
 AND4_X1 _28371_ (.A1(_04703_),
    .A2(_04906_),
    .A3(_04903_),
    .A4(_04907_),
    .ZN(_04961_));
 NOR4_X2 _28372_ (.A1(_04662_),
    .A2(_04717_),
    .A3(_04907_),
    .A4(_04895_),
    .ZN(_04962_));
 NAND2_X1 _28373_ (.A1(_04696_),
    .A2(_04698_),
    .ZN(_04963_));
 NAND2_X1 _28374_ (.A1(_04699_),
    .A2(_04702_),
    .ZN(_04964_));
 OAI33_X1 _28375_ (.A1(_04650_),
    .A2(_04658_),
    .A3(_04660_),
    .B1(_04963_),
    .B2(_04964_),
    .B3(_04955_),
    .ZN(_04965_));
 AOI211_X2 _28376_ (.A(_04961_),
    .B(_04962_),
    .C1(_04906_),
    .C2(_04965_),
    .ZN(_04966_));
 AOI221_X2 _28377_ (.A(_04941_),
    .B1(_04948_),
    .B2(_04950_),
    .C1(_04960_),
    .C2(_04966_),
    .ZN(_04967_));
 NAND2_X2 _28378_ (.A1(_04924_),
    .A2(_04929_),
    .ZN(_04968_));
 OAI21_X4 _28379_ (.A(_04940_),
    .B1(_04967_),
    .B2(_04968_),
    .ZN(_04969_));
 CLKBUF_X3 _28380_ (.A(_14179_),
    .Z(_04970_));
 INV_X1 _28381_ (.A(_04970_),
    .ZN(_04971_));
 XNOR2_X2 _28382_ (.A(_04837_),
    .B(_04804_),
    .ZN(_04972_));
 OR3_X1 _28383_ (.A1(_04863_),
    .A2(_04868_),
    .A3(_04891_),
    .ZN(_04973_));
 AOI21_X1 _28384_ (.A(_04973_),
    .B1(_04953_),
    .B2(_04959_),
    .ZN(_04974_));
 INV_X1 _28385_ (.A(_04880_),
    .ZN(_04975_));
 BUF_X2 _28386_ (.A(_04868_),
    .Z(_04976_));
 NOR2_X1 _28387_ (.A1(_04949_),
    .A2(_04976_),
    .ZN(_04977_));
 AOI221_X2 _28388_ (.A(_04972_),
    .B1(_04974_),
    .B2(_04966_),
    .C1(_04975_),
    .C2(_04977_),
    .ZN(_04978_));
 NOR3_X2 _28389_ (.A1(_04971_),
    .A2(_04893_),
    .A3(_04978_),
    .ZN(_04979_));
 NOR3_X4 _28390_ (.A1(_04661_),
    .A2(_04717_),
    .A3(_04836_),
    .ZN(_04980_));
 XNOR2_X2 _28391_ (.A(_04980_),
    .B(_04804_),
    .ZN(_04981_));
 NOR3_X1 _28392_ (.A1(_04949_),
    .A2(_04976_),
    .A3(_04891_),
    .ZN(_04982_));
 OAI21_X1 _28393_ (.A(_04982_),
    .B1(_04896_),
    .B2(_04904_),
    .ZN(_04983_));
 OAI221_X2 _28394_ (.A(_04981_),
    .B1(_04983_),
    .B2(_04912_),
    .C1(_04880_),
    .C2(_04869_),
    .ZN(_04984_));
 NAND3_X1 _28395_ (.A1(_04703_),
    .A2(_04903_),
    .A3(_04907_),
    .ZN(_04985_));
 NAND2_X2 _28396_ (.A1(_04911_),
    .A2(_04985_),
    .ZN(_04986_));
 XNOR2_X2 _28397_ (.A(_04781_),
    .B(_04986_),
    .ZN(_04987_));
 AOI21_X1 _28398_ (.A(_04984_),
    .B1(_04987_),
    .B2(_04970_),
    .ZN(_04988_));
 BUF_X1 _28399_ (.A(_22250_),
    .Z(_04989_));
 NOR2_X1 _28400_ (.A1(_04989_),
    .A2(_04893_),
    .ZN(_04990_));
 NOR2_X1 _28401_ (.A1(_04837_),
    .A2(_04934_),
    .ZN(_04991_));
 NOR2_X1 _28402_ (.A1(_04980_),
    .A2(_04935_),
    .ZN(_04992_));
 OAI33_X1 _28403_ (.A1(_04969_),
    .A2(_04979_),
    .A3(_04988_),
    .B1(_04990_),
    .B2(_04991_),
    .B3(_04992_),
    .ZN(_04993_));
 CLKBUF_X3 _28404_ (.A(_04970_),
    .Z(_04994_));
 OAI21_X1 _28405_ (.A(_04994_),
    .B1(_04978_),
    .B2(_04987_),
    .ZN(_04995_));
 BUF_X4 _28406_ (.A(_04936_),
    .Z(_04996_));
 OAI21_X1 _28407_ (.A(_04996_),
    .B1(_04987_),
    .B2(_04989_),
    .ZN(_04997_));
 NAND2_X1 _28408_ (.A1(_04989_),
    .A2(_04996_),
    .ZN(_04998_));
 AOI21_X1 _28409_ (.A(_04998_),
    .B1(_04945_),
    .B2(_04893_),
    .ZN(_04999_));
 OAI22_X1 _28410_ (.A1(_04969_),
    .A2(_04995_),
    .B1(_04997_),
    .B2(_04999_),
    .ZN(_05000_));
 AND2_X1 _28411_ (.A1(_04993_),
    .A2(_05000_),
    .ZN(_22256_));
 BUF_X4 _28412_ (.A(_04585_),
    .Z(_05001_));
 NOR2_X1 _28413_ (.A1(\g_reduce0[6].adder.x[0] ),
    .A2(_05001_),
    .ZN(_05002_));
 NOR4_X4 _28414_ (.A1(_04581_),
    .A2(_04582_),
    .A3(_04583_),
    .A4(_04584_),
    .ZN(_05003_));
 AOI21_X1 _28415_ (.A(_05003_),
    .B1(_04589_),
    .B2(\g_reduce0[4].adder.x[0] ),
    .ZN(_05004_));
 INV_X2 _28416_ (.A(_04589_),
    .ZN(_05005_));
 OAI21_X1 _28417_ (.A(_04997_),
    .B1(_04995_),
    .B2(_04969_),
    .ZN(_05006_));
 NAND3_X1 _28418_ (.A1(_04920_),
    .A2(_04921_),
    .A3(_04923_),
    .ZN(_05007_));
 NOR2_X1 _28419_ (.A1(_05007_),
    .A2(_04996_),
    .ZN(_05008_));
 NAND2_X1 _28420_ (.A1(_04948_),
    .A2(_04950_),
    .ZN(_05009_));
 NOR2_X1 _28421_ (.A1(_04949_),
    .A2(_04951_),
    .ZN(_05010_));
 OAI21_X1 _28422_ (.A(_05010_),
    .B1(_04896_),
    .B2(_04904_),
    .ZN(_05011_));
 OAI211_X2 _28423_ (.A(_04919_),
    .B(_05009_),
    .C1(_05011_),
    .C2(_04912_),
    .ZN(_05012_));
 AOI21_X4 _28424_ (.A(_04872_),
    .B1(_05008_),
    .B2(_05012_),
    .ZN(_22279_));
 AND3_X1 _28425_ (.A1(_22252_),
    .A2(_22275_),
    .A3(_22279_),
    .ZN(_05013_));
 OAI221_X1 _28426_ (.A(_05006_),
    .B1(_05013_),
    .B2(_04996_),
    .C1(_04998_),
    .C2(_04893_),
    .ZN(_05014_));
 OAI21_X1 _28427_ (.A(_04993_),
    .B1(_04998_),
    .B2(_04945_),
    .ZN(_05015_));
 AOI21_X1 _28428_ (.A(_22256_),
    .B1(_05014_),
    .B2(_05015_),
    .ZN(_05016_));
 CLKBUF_X3 _28429_ (.A(_04989_),
    .Z(_05017_));
 AOI21_X4 _28430_ (.A(_04833_),
    .B1(_04980_),
    .B2(_04820_),
    .ZN(_05018_));
 BUF_X4 _28431_ (.A(_05018_),
    .Z(_05019_));
 CLKBUF_X3 _28432_ (.A(_04971_),
    .Z(_14174_));
 AND2_X1 _28433_ (.A1(_22245_),
    .A2(_04785_),
    .ZN(_05020_));
 AOI21_X1 _28434_ (.A(_05020_),
    .B1(_04781_),
    .B2(_22247_),
    .ZN(_05021_));
 NOR2_X1 _28435_ (.A1(_05021_),
    .A2(_04950_),
    .ZN(_05022_));
 NOR2_X1 _28436_ (.A1(_04949_),
    .A2(_04891_),
    .ZN(_05023_));
 OAI21_X1 _28437_ (.A(_05023_),
    .B1(_04896_),
    .B2(_04904_),
    .ZN(_05024_));
 OAI211_X2 _28438_ (.A(_04929_),
    .B(_05022_),
    .C1(_05024_),
    .C2(_04912_),
    .ZN(_05025_));
 OR2_X2 _28439_ (.A1(_04869_),
    .A2(_04872_),
    .ZN(_05026_));
 NOR2_X2 _28440_ (.A1(_05026_),
    .A2(_04886_),
    .ZN(_05027_));
 NOR2_X1 _28441_ (.A1(_04921_),
    .A2(_05021_),
    .ZN(_05028_));
 MUX2_X1 _28442_ (.A(_04945_),
    .B(_05028_),
    .S(_04981_),
    .Z(_05029_));
 AOI22_X4 _28443_ (.A1(_04913_),
    .A2(_05027_),
    .B1(_05029_),
    .B2(_05019_),
    .ZN(_05030_));
 NAND2_X1 _28444_ (.A1(_05025_),
    .A2(_05030_),
    .ZN(_05031_));
 NAND3_X1 _28445_ (.A1(_14174_),
    .A2(_04940_),
    .A3(_05031_),
    .ZN(_05032_));
 OAI22_X1 _28446_ (.A1(_05017_),
    .A2(_05019_),
    .B1(_22279_),
    .B2(_05032_),
    .ZN(_05033_));
 AOI21_X1 _28447_ (.A(_04936_),
    .B1(_04924_),
    .B2(_04941_),
    .ZN(_05034_));
 NOR2_X1 _28448_ (.A1(_04904_),
    .A2(_04896_),
    .ZN(_05035_));
 OR4_X1 _28449_ (.A1(_04912_),
    .A2(_05035_),
    .A3(_05007_),
    .A4(_04951_),
    .ZN(_05036_));
 AND2_X1 _28450_ (.A1(_05034_),
    .A2(_05036_),
    .ZN(_05037_));
 INV_X1 _28451_ (.A(_04875_),
    .ZN(_05038_));
 NOR3_X1 _28452_ (.A1(_04804_),
    .A2(_05038_),
    .A3(_04921_),
    .ZN(_05039_));
 AOI22_X2 _28453_ (.A1(_04922_),
    .A2(_04875_),
    .B1(_05039_),
    .B2(_04836_),
    .ZN(_05040_));
 NOR2_X1 _28454_ (.A1(_04920_),
    .A2(_04976_),
    .ZN(_05041_));
 NOR2_X1 _28455_ (.A1(_04972_),
    .A2(_05041_),
    .ZN(_05042_));
 NOR3_X1 _28456_ (.A1(_04719_),
    .A2(_04836_),
    .A3(_04834_),
    .ZN(_05043_));
 AOI21_X1 _28457_ (.A(_05043_),
    .B1(_04834_),
    .B2(_04719_),
    .ZN(_05044_));
 NAND2_X1 _28458_ (.A1(_04875_),
    .A2(_04976_),
    .ZN(_05045_));
 OAI221_X2 _28459_ (.A(_05040_),
    .B1(_05042_),
    .B2(_04847_),
    .C1(_05044_),
    .C2(_05045_),
    .ZN(_05046_));
 NOR2_X1 _28460_ (.A1(_04971_),
    .A2(_04872_),
    .ZN(_05047_));
 NAND3_X1 _28461_ (.A1(_04938_),
    .A2(_05046_),
    .A3(_05047_),
    .ZN(_05048_));
 INV_X1 _28462_ (.A(_04920_),
    .ZN(_05049_));
 NAND4_X1 _28463_ (.A1(_14174_),
    .A2(_05049_),
    .A3(_04976_),
    .A4(_22275_),
    .ZN(_05050_));
 NOR3_X1 _28464_ (.A1(_04804_),
    .A2(_04921_),
    .A3(_04918_),
    .ZN(_05051_));
 NOR3_X1 _28465_ (.A1(_04834_),
    .A2(_04921_),
    .A3(_04918_),
    .ZN(_05052_));
 MUX2_X1 _28466_ (.A(_05051_),
    .B(_05052_),
    .S(_04980_),
    .Z(_05053_));
 OAI21_X1 _28467_ (.A(_04834_),
    .B1(_04949_),
    .B2(_04976_),
    .ZN(_05054_));
 OAI21_X1 _28468_ (.A(_04804_),
    .B1(_04949_),
    .B2(_04976_),
    .ZN(_05055_));
 MUX2_X1 _28469_ (.A(_05054_),
    .B(_05055_),
    .S(_04980_),
    .Z(_05056_));
 NOR2_X1 _28470_ (.A1(_04916_),
    .A2(_04872_),
    .ZN(_05057_));
 AND2_X1 _28471_ (.A1(_04949_),
    .A2(_04879_),
    .ZN(_05058_));
 AOI222_X2 _28472_ (.A1(_05018_),
    .A2(_05053_),
    .B1(_05056_),
    .B2(_05057_),
    .C1(_05058_),
    .C2(_04929_),
    .ZN(_05059_));
 OR3_X1 _28473_ (.A1(_04994_),
    .A2(_22275_),
    .A3(_05059_),
    .ZN(_05060_));
 NAND3_X1 _28474_ (.A1(_05048_),
    .A2(_05050_),
    .A3(_05060_),
    .ZN(_05061_));
 AND2_X1 _28475_ (.A1(_05037_),
    .A2(_05061_),
    .ZN(_05062_));
 OAI21_X1 _28476_ (.A(_04890_),
    .B1(_04880_),
    .B2(_04949_),
    .ZN(_05063_));
 OR2_X1 _28477_ (.A1(_04863_),
    .A2(_04891_),
    .ZN(_05064_));
 AOI21_X1 _28478_ (.A(_05064_),
    .B1(_04953_),
    .B2(_04959_),
    .ZN(_05065_));
 AOI211_X2 _28479_ (.A(_04936_),
    .B(_05063_),
    .C1(_05065_),
    .C2(_04966_),
    .ZN(_05066_));
 NOR2_X1 _28480_ (.A1(_05026_),
    .A2(_04885_),
    .ZN(_05067_));
 NOR2_X1 _28481_ (.A1(_04921_),
    .A2(_04917_),
    .ZN(_05068_));
 MUX2_X1 _28482_ (.A(_04943_),
    .B(_05068_),
    .S(_04981_),
    .Z(_05069_));
 AOI221_X2 _28483_ (.A(_05066_),
    .B1(_05067_),
    .B2(_04913_),
    .C1(_05018_),
    .C2(_05069_),
    .ZN(_05070_));
 NAND2_X1 _28484_ (.A1(_05019_),
    .A2(_04978_),
    .ZN(_05071_));
 AOI211_X4 _28485_ (.A(_04930_),
    .B(_04937_),
    .C1(_04987_),
    .C2(_05018_),
    .ZN(_05072_));
 AOI22_X4 _28486_ (.A1(_22275_),
    .A2(_05070_),
    .B1(_05071_),
    .B2(_05072_),
    .ZN(_05073_));
 NAND2_X2 _28487_ (.A1(_04970_),
    .A2(_05019_),
    .ZN(_05074_));
 NOR4_X2 _28488_ (.A1(_04972_),
    .A2(_04968_),
    .A3(_04967_),
    .A4(_05074_),
    .ZN(_05075_));
 AOI211_X2 _28489_ (.A(_05033_),
    .B(_05062_),
    .C1(_05073_),
    .C2(_05075_),
    .ZN(_05076_));
 NAND2_X1 _28490_ (.A1(_04938_),
    .A2(_05037_),
    .ZN(_05077_));
 MUX2_X1 _28491_ (.A(_05059_),
    .B(_05070_),
    .S(_14174_),
    .Z(_05078_));
 OR2_X1 _28492_ (.A1(_05077_),
    .A2(_05078_),
    .ZN(_05079_));
 AOI21_X1 _28493_ (.A(_04921_),
    .B1(_04981_),
    .B2(_04920_),
    .ZN(_05080_));
 MUX2_X1 _28494_ (.A(_05046_),
    .B(_05080_),
    .S(_04994_),
    .Z(_05081_));
 MUX2_X1 _28495_ (.A(_04976_),
    .B(_04972_),
    .S(_05017_),
    .Z(_05082_));
 AOI22_X2 _28496_ (.A1(_04940_),
    .A2(_05081_),
    .B1(_05082_),
    .B2(_04996_),
    .ZN(_05083_));
 CLKBUF_X3 _28497_ (.A(_04929_),
    .Z(_05084_));
 NAND2_X1 _28498_ (.A1(_05084_),
    .A2(_04939_),
    .ZN(_05085_));
 XNOR2_X2 _28499_ (.A(_04785_),
    .B(_04986_),
    .ZN(_05086_));
 AOI21_X1 _28500_ (.A(_04872_),
    .B1(_04984_),
    .B2(_05086_),
    .ZN(_05087_));
 NOR2_X1 _28501_ (.A1(_04994_),
    .A2(_05087_),
    .ZN(_05088_));
 AND3_X1 _28502_ (.A1(_04994_),
    .A2(_05025_),
    .A3(_05030_),
    .ZN(_05089_));
 OR4_X1 _28503_ (.A1(_05085_),
    .A2(_22279_),
    .A3(_05088_),
    .A4(_05089_),
    .ZN(_05090_));
 NAND3_X2 _28504_ (.A1(_05079_),
    .A2(_05083_),
    .A3(_05090_),
    .ZN(_05091_));
 MUX2_X1 _28505_ (.A(_05049_),
    .B(_04976_),
    .S(_05017_),
    .Z(_05092_));
 NOR3_X2 _28506_ (.A1(_04922_),
    .A2(_04875_),
    .A3(_04948_),
    .ZN(_05093_));
 NAND2_X1 _28507_ (.A1(_04920_),
    .A2(_04921_),
    .ZN(_05094_));
 OAI21_X4 _28508_ (.A(_04929_),
    .B1(_05093_),
    .B2(_05094_),
    .ZN(_22248_));
 NAND3_X2 _28509_ (.A1(_04914_),
    .A2(_04919_),
    .A3(_22248_),
    .ZN(_05095_));
 OAI22_X4 _28510_ (.A1(_04914_),
    .A2(_04919_),
    .B1(_05095_),
    .B2(_22249_),
    .ZN(_05096_));
 AOI221_X2 _28511_ (.A(_04838_),
    .B1(_04873_),
    .B2(_04913_),
    .C1(_04987_),
    .C2(_05047_),
    .ZN(_05097_));
 NOR3_X2 _28512_ (.A1(_04968_),
    .A2(_04979_),
    .A3(_05097_),
    .ZN(_05098_));
 AOI22_X4 _28513_ (.A1(_04996_),
    .A2(_05092_),
    .B1(_05096_),
    .B2(_05098_),
    .ZN(_05099_));
 NAND2_X1 _28514_ (.A1(_05034_),
    .A2(_05036_),
    .ZN(_05100_));
 OAI21_X1 _28515_ (.A(_04933_),
    .B1(_04803_),
    .B2(_04782_),
    .ZN(_05101_));
 NOR4_X1 _28516_ (.A1(_04662_),
    .A2(_04717_),
    .A3(_04836_),
    .A4(_05101_),
    .ZN(_05102_));
 AOI21_X1 _28517_ (.A(_05102_),
    .B1(_04835_),
    .B2(_04837_),
    .ZN(_05103_));
 NAND2_X1 _28518_ (.A1(_05103_),
    .A2(_05026_),
    .ZN(_05104_));
 NOR2_X1 _28519_ (.A1(_04838_),
    .A2(_04885_),
    .ZN(_05105_));
 NAND2_X1 _28520_ (.A1(_04873_),
    .A2(_04975_),
    .ZN(_05106_));
 AOI221_X2 _28521_ (.A(_14174_),
    .B1(_04879_),
    .B2(_05104_),
    .C1(_05105_),
    .C2(_05106_),
    .ZN(_05107_));
 NOR3_X1 _28522_ (.A1(_22275_),
    .A2(_05100_),
    .A3(_05107_),
    .ZN(_05108_));
 MUX2_X1 _28523_ (.A(_04890_),
    .B(_04945_),
    .S(_22249_),
    .Z(_05109_));
 OAI21_X2 _28524_ (.A(_05108_),
    .B1(_05109_),
    .B2(_04994_),
    .ZN(_05110_));
 MUX2_X1 _28525_ (.A(_05049_),
    .B(_04922_),
    .S(_04981_),
    .Z(_05111_));
 OR3_X1 _28526_ (.A1(_14174_),
    .A2(_05041_),
    .A3(_05111_),
    .ZN(_05112_));
 AOI211_X2 _28527_ (.A(_04838_),
    .B(_04942_),
    .C1(_04873_),
    .C2(_04913_),
    .ZN(_05113_));
 AOI21_X2 _28528_ (.A(_05113_),
    .B1(_22251_),
    .B2(_05038_),
    .ZN(_05114_));
 OAI21_X2 _28529_ (.A(_05112_),
    .B1(_05114_),
    .B2(_04994_),
    .ZN(_05115_));
 OAI211_X4 _28530_ (.A(_05099_),
    .B(_05110_),
    .C1(_05115_),
    .C2(_04969_),
    .ZN(_05116_));
 INV_X2 _28531_ (.A(_04989_),
    .ZN(_05117_));
 MUX2_X1 _28532_ (.A(_05019_),
    .B(_04981_),
    .S(_05117_),
    .Z(_05118_));
 NOR3_X1 _28533_ (.A1(_04970_),
    .A2(_05041_),
    .A3(_05111_),
    .ZN(_05119_));
 NOR3_X1 _28534_ (.A1(_04971_),
    .A2(_04976_),
    .A3(_04972_),
    .ZN(_05120_));
 NOR4_X1 _28535_ (.A1(_04872_),
    .A2(_04938_),
    .A3(_05119_),
    .A4(_05120_),
    .ZN(_05121_));
 NAND2_X1 _28536_ (.A1(_04879_),
    .A2(_05104_),
    .ZN(_05122_));
 NAND2_X1 _28537_ (.A1(_05105_),
    .A2(_05106_),
    .ZN(_05123_));
 AOI21_X1 _28538_ (.A(_04994_),
    .B1(_05122_),
    .B2(_05123_),
    .ZN(_05124_));
 AOI21_X1 _28539_ (.A(_05121_),
    .B1(_05124_),
    .B2(_04938_),
    .ZN(_05125_));
 NAND2_X1 _28540_ (.A1(_22279_),
    .A2(_05118_),
    .ZN(_05126_));
 NOR2_X1 _28541_ (.A1(_14174_),
    .A2(_22275_),
    .ZN(_05127_));
 AOI21_X1 _28542_ (.A(_05126_),
    .B1(_05127_),
    .B2(_05114_),
    .ZN(_05128_));
 INV_X1 _28543_ (.A(_05118_),
    .ZN(_05129_));
 NOR2_X1 _28544_ (.A1(_22279_),
    .A2(_05129_),
    .ZN(_05130_));
 NOR2_X1 _28545_ (.A1(_04917_),
    .A2(_05074_),
    .ZN(_05131_));
 NOR2_X1 _28546_ (.A1(_04886_),
    .A2(_05074_),
    .ZN(_05132_));
 MUX2_X1 _28547_ (.A(_05131_),
    .B(_05132_),
    .S(_22249_),
    .Z(_05133_));
 NOR2_X1 _28548_ (.A1(_14179_),
    .A2(_04872_),
    .ZN(_05134_));
 OAI21_X1 _28549_ (.A(_05134_),
    .B1(_04981_),
    .B2(_04893_),
    .ZN(_05135_));
 NOR2_X1 _28550_ (.A1(_05026_),
    .A2(_04893_),
    .ZN(_05136_));
 AOI221_X2 _28551_ (.A(_05135_),
    .B1(_05086_),
    .B2(_04978_),
    .C1(_04913_),
    .C2(_05136_),
    .ZN(_05137_));
 OR2_X1 _28552_ (.A1(_04938_),
    .A2(_05137_),
    .ZN(_05138_));
 OAI22_X1 _28553_ (.A1(_22252_),
    .A2(_22275_),
    .B1(_05133_),
    .B2(_05138_),
    .ZN(_05139_));
 AOI222_X4 _28554_ (.A1(_04996_),
    .A2(_05118_),
    .B1(_05125_),
    .B2(_05128_),
    .C1(_05130_),
    .C2(_05139_),
    .ZN(_05140_));
 NAND3_X1 _28555_ (.A1(_05091_),
    .A2(_05116_),
    .A3(_05140_),
    .ZN(_05141_));
 AOI21_X1 _28556_ (.A(_04994_),
    .B1(_04890_),
    .B2(_22251_),
    .ZN(_05142_));
 OR3_X1 _28557_ (.A1(_04969_),
    .A2(_05107_),
    .A3(_05142_),
    .ZN(_05143_));
 NOR4_X1 _28558_ (.A1(_22275_),
    .A2(_05100_),
    .A3(_04979_),
    .A4(_05097_),
    .ZN(_05144_));
 MUX2_X1 _28559_ (.A(_04942_),
    .B(_04879_),
    .S(_05117_),
    .Z(_05145_));
 AOI21_X1 _28560_ (.A(_05144_),
    .B1(_05145_),
    .B2(_04996_),
    .ZN(_05146_));
 NOR2_X1 _28561_ (.A1(_04970_),
    .A2(_04969_),
    .ZN(_05147_));
 NAND4_X1 _28562_ (.A1(_05019_),
    .A2(_04945_),
    .A3(_22249_),
    .A4(_05147_),
    .ZN(_05148_));
 NAND3_X2 _28563_ (.A1(_05143_),
    .A2(_05146_),
    .A3(_05148_),
    .ZN(_05149_));
 NOR2_X1 _28564_ (.A1(_04879_),
    .A2(_04998_),
    .ZN(_05150_));
 AOI21_X1 _28565_ (.A(_04929_),
    .B1(_04885_),
    .B2(_05117_),
    .ZN(_05151_));
 AND3_X1 _28566_ (.A1(_04970_),
    .A2(_05034_),
    .A3(_05036_),
    .ZN(_05152_));
 AOI221_X2 _28567_ (.A(_05151_),
    .B1(_05147_),
    .B2(_05031_),
    .C1(_05152_),
    .C2(_05073_),
    .ZN(_05153_));
 MUX2_X1 _28568_ (.A(_04890_),
    .B(_04943_),
    .S(_05017_),
    .Z(_05154_));
 NAND2_X1 _28569_ (.A1(_04996_),
    .A2(_05154_),
    .ZN(_05155_));
 INV_X1 _28570_ (.A(_22252_),
    .ZN(_05156_));
 AOI21_X1 _28571_ (.A(_05100_),
    .B1(_04938_),
    .B2(_05156_),
    .ZN(_05157_));
 OAI21_X1 _28572_ (.A(_05157_),
    .B1(_05138_),
    .B2(_05133_),
    .ZN(_05158_));
 AOI211_X4 _28573_ (.A(_05150_),
    .B(_05153_),
    .C1(_05155_),
    .C2(_05158_),
    .ZN(_05159_));
 NAND2_X1 _28574_ (.A1(_05017_),
    .A2(_04920_),
    .ZN(_05160_));
 OAI221_X2 _28575_ (.A(_05160_),
    .B1(_04972_),
    .B2(_04872_),
    .C1(_05017_),
    .C2(_04922_),
    .ZN(_05161_));
 AND2_X1 _28576_ (.A1(_05025_),
    .A2(_05030_),
    .ZN(_05162_));
 MUX2_X1 _28577_ (.A(_05162_),
    .B(_05070_),
    .S(_04994_),
    .Z(_05163_));
 NAND2_X1 _28578_ (.A1(_14174_),
    .A2(_05059_),
    .ZN(_05164_));
 MUX2_X1 _28579_ (.A(_05087_),
    .B(_05046_),
    .S(_22279_),
    .Z(_05165_));
 OAI21_X1 _28580_ (.A(_05164_),
    .B1(_05165_),
    .B2(_14174_),
    .ZN(_05166_));
 OAI221_X2 _28581_ (.A(_05161_),
    .B1(_05163_),
    .B2(_05077_),
    .C1(_05166_),
    .C2(_05085_),
    .ZN(_05167_));
 AOI211_X2 _28582_ (.A(_05074_),
    .B(_05113_),
    .C1(_05038_),
    .C2(_22251_),
    .ZN(_05168_));
 NAND2_X1 _28583_ (.A1(_14174_),
    .A2(_05019_),
    .ZN(_05169_));
 AOI21_X1 _28584_ (.A(_05169_),
    .B1(_05122_),
    .B2(_05123_),
    .ZN(_05170_));
 OAI33_X1 _28585_ (.A1(_05133_),
    .A2(_05137_),
    .A3(_05077_),
    .B1(_05168_),
    .B2(_05170_),
    .B3(_04969_),
    .ZN(_05171_));
 MUX2_X1 _28586_ (.A(_04922_),
    .B(_04875_),
    .S(_05117_),
    .Z(_05172_));
 OAI21_X1 _28587_ (.A(_05084_),
    .B1(_04938_),
    .B2(_05156_),
    .ZN(_05173_));
 OAI22_X2 _28588_ (.A1(_05084_),
    .A2(_05172_),
    .B1(_05173_),
    .B2(_22279_),
    .ZN(_05174_));
 NOR2_X1 _28589_ (.A1(_05117_),
    .A2(_04875_),
    .ZN(_05175_));
 AOI221_X2 _28590_ (.A(_05175_),
    .B1(_04981_),
    .B2(_05019_),
    .C1(_05117_),
    .C2(_04916_),
    .ZN(_05176_));
 NAND3_X1 _28591_ (.A1(_04938_),
    .A2(_05025_),
    .A3(_05030_),
    .ZN(_05177_));
 OAI21_X1 _28592_ (.A(_05059_),
    .B1(_04937_),
    .B2(_04930_),
    .ZN(_05178_));
 AND2_X1 _28593_ (.A1(_05152_),
    .A2(_05178_),
    .ZN(_05179_));
 NOR2_X1 _28594_ (.A1(_04970_),
    .A2(_05100_),
    .ZN(_05180_));
 AOI221_X2 _28595_ (.A(_05176_),
    .B1(_05177_),
    .B2(_05179_),
    .C1(_05073_),
    .C2(_05180_),
    .ZN(_05181_));
 MUX2_X1 _28596_ (.A(_04890_),
    .B(_04945_),
    .S(_05117_),
    .Z(_05182_));
 NAND2_X1 _28597_ (.A1(_04936_),
    .A2(_05182_),
    .ZN(_05183_));
 AOI21_X1 _28598_ (.A(_04970_),
    .B1(_04996_),
    .B2(_05182_),
    .ZN(_05184_));
 OAI21_X1 _28599_ (.A(_05019_),
    .B1(_04978_),
    .B2(_04987_),
    .ZN(_05185_));
 AND3_X1 _28600_ (.A1(_04970_),
    .A2(_05025_),
    .A3(_05183_),
    .ZN(_05186_));
 AOI222_X2 _28601_ (.A1(_04969_),
    .A2(_05183_),
    .B1(_05184_),
    .B2(_05185_),
    .C1(_05186_),
    .C2(_05030_),
    .ZN(_22257_));
 NAND3_X1 _28602_ (.A1(_04993_),
    .A2(_05000_),
    .A3(_22257_),
    .ZN(_05187_));
 NOR4_X2 _28603_ (.A1(_05171_),
    .A2(_05174_),
    .A3(_05181_),
    .A4(_05187_),
    .ZN(_05188_));
 NAND4_X2 _28604_ (.A1(_05149_),
    .A2(_05159_),
    .A3(_05167_),
    .A4(_05188_),
    .ZN(_05189_));
 NOR2_X1 _28605_ (.A1(_05141_),
    .A2(_05189_),
    .ZN(_05190_));
 XNOR2_X2 _28606_ (.A(_05076_),
    .B(_05190_),
    .ZN(_22262_));
 MUX2_X1 _28607_ (.A(_05016_),
    .B(_22259_),
    .S(_22262_),
    .Z(_05191_));
 NAND2_X1 _28608_ (.A1(_05005_),
    .A2(_05191_),
    .ZN(_05192_));
 AOI21_X1 _28609_ (.A(_05002_),
    .B1(_05004_),
    .B2(_05192_),
    .ZN(_00144_));
 NOR2_X4 _28610_ (.A1(_05003_),
    .A2(_04589_),
    .ZN(_05193_));
 NAND2_X1 _28611_ (.A1(_22259_),
    .A2(_05193_),
    .ZN(_05194_));
 NAND2_X1 _28612_ (.A1(_05155_),
    .A2(_05158_),
    .ZN(_05195_));
 XOR2_X1 _28613_ (.A(_22258_),
    .B(_05195_),
    .Z(_05196_));
 NAND2_X1 _28614_ (.A1(_05193_),
    .A2(_05196_),
    .ZN(_05197_));
 MUX2_X1 _28615_ (.A(_05194_),
    .B(_05197_),
    .S(_22262_),
    .Z(_05198_));
 NOR2_X2 _28616_ (.A1(_05003_),
    .A2(_05005_),
    .ZN(_05199_));
 AOI22_X2 _28617_ (.A1(\g_reduce0[6].adder.x[1] ),
    .A2(_05003_),
    .B1(_05199_),
    .B2(\g_reduce0[4].adder.x[1] ),
    .ZN(_05200_));
 NAND2_X1 _28618_ (.A1(_05198_),
    .A2(_05200_),
    .ZN(_00151_));
 OR2_X1 _28619_ (.A1(_22262_),
    .A2(_05197_),
    .ZN(_05201_));
 NOR2_X1 _28620_ (.A1(_05150_),
    .A2(_05153_),
    .ZN(_05202_));
 INV_X1 _28621_ (.A(_05187_),
    .ZN(_05203_));
 NAND2_X1 _28622_ (.A1(_05195_),
    .A2(_05203_),
    .ZN(_05204_));
 XNOR2_X1 _28623_ (.A(_05202_),
    .B(_05204_),
    .ZN(_05205_));
 NAND3_X1 _28624_ (.A1(_22262_),
    .A2(_05193_),
    .A3(_05205_),
    .ZN(_05206_));
 AOI22_X2 _28625_ (.A1(\g_reduce0[6].adder.x[2] ),
    .A2(_05003_),
    .B1(_05199_),
    .B2(\g_reduce0[4].adder.x[2] ),
    .ZN(_05207_));
 NAND3_X1 _28626_ (.A1(_05201_),
    .A2(_05206_),
    .A3(_05207_),
    .ZN(_00152_));
 NAND2_X2 _28627_ (.A1(_04585_),
    .A2(_04589_),
    .ZN(_05208_));
 OAI22_X2 _28628_ (.A1(\g_reduce0[6].adder.x[3] ),
    .A2(_05001_),
    .B1(_05208_),
    .B2(\g_reduce0[4].adder.x[3] ),
    .ZN(_05209_));
 NAND2_X1 _28629_ (.A1(_22258_),
    .A2(_05159_),
    .ZN(_05210_));
 XOR2_X1 _28630_ (.A(_05149_),
    .B(_05210_),
    .Z(_05211_));
 NAND2_X1 _28631_ (.A1(_22262_),
    .A2(_05211_),
    .ZN(_05212_));
 OAI21_X1 _28632_ (.A(_05212_),
    .B1(_05205_),
    .B2(_22262_),
    .ZN(_05213_));
 AOI21_X1 _28633_ (.A(_05209_),
    .B1(_05213_),
    .B2(_05193_),
    .ZN(_00153_));
 AOI22_X2 _28634_ (.A1(\g_reduce0[6].adder.x[4] ),
    .A2(_05003_),
    .B1(_05199_),
    .B2(\g_reduce0[4].adder.x[4] ),
    .ZN(_05214_));
 NAND2_X1 _28635_ (.A1(_05073_),
    .A2(_05180_),
    .ZN(_05215_));
 AOI21_X1 _28636_ (.A(_05176_),
    .B1(_05177_),
    .B2(_05179_),
    .ZN(_05216_));
 NAND2_X1 _28637_ (.A1(_05215_),
    .A2(_05216_),
    .ZN(_05217_));
 AND3_X1 _28638_ (.A1(_05149_),
    .A2(_05159_),
    .A3(_05203_),
    .ZN(_05218_));
 XNOR2_X1 _28639_ (.A(_05217_),
    .B(_05218_),
    .ZN(_05219_));
 MUX2_X1 _28640_ (.A(_05211_),
    .B(_05219_),
    .S(_22262_),
    .Z(_05220_));
 NAND2_X1 _28641_ (.A1(_04585_),
    .A2(_05005_),
    .ZN(_05221_));
 OAI21_X1 _28642_ (.A(_05214_),
    .B1(_05220_),
    .B2(_05221_),
    .ZN(_00154_));
 OAI22_X2 _28643_ (.A1(\g_reduce0[6].adder.x[5] ),
    .A2(_05001_),
    .B1(_05208_),
    .B2(\g_reduce0[4].adder.x[5] ),
    .ZN(_05222_));
 NOR2_X1 _28644_ (.A1(_05171_),
    .A2(_05174_),
    .ZN(_05223_));
 AND4_X1 _28645_ (.A1(_22258_),
    .A2(_05149_),
    .A3(_05159_),
    .A4(_05217_),
    .ZN(_05224_));
 XNOR2_X1 _28646_ (.A(_05223_),
    .B(_05224_),
    .ZN(_05225_));
 MUX2_X1 _28647_ (.A(_05219_),
    .B(_05225_),
    .S(_22262_),
    .Z(_05226_));
 AOI21_X1 _28648_ (.A(_05222_),
    .B1(_05226_),
    .B2(_05193_),
    .ZN(_00155_));
 OAI22_X2 _28649_ (.A1(\g_reduce0[6].adder.x[6] ),
    .A2(_05001_),
    .B1(_05208_),
    .B2(\g_reduce0[4].adder.x[6] ),
    .ZN(_05227_));
 BUF_X2 _28650_ (.A(_05076_),
    .Z(_05228_));
 AND3_X1 _28651_ (.A1(_05149_),
    .A2(_05159_),
    .A3(_05188_),
    .ZN(_05229_));
 XNOR2_X1 _28652_ (.A(_05167_),
    .B(_05229_),
    .ZN(_05230_));
 OR3_X1 _28653_ (.A1(_05141_),
    .A2(_05189_),
    .A3(_05225_),
    .ZN(_05231_));
 AOI21_X1 _28654_ (.A(_05228_),
    .B1(_05230_),
    .B2(_05231_),
    .ZN(_05232_));
 NOR2_X1 _28655_ (.A1(_05190_),
    .A2(_05225_),
    .ZN(_05233_));
 AOI21_X1 _28656_ (.A(_05232_),
    .B1(_05233_),
    .B2(_05228_),
    .ZN(_05234_));
 AOI21_X1 _28657_ (.A(_05227_),
    .B1(_05234_),
    .B2(_05193_),
    .ZN(_00156_));
 AOI22_X2 _28658_ (.A1(\g_reduce0[6].adder.x[7] ),
    .A2(_05003_),
    .B1(_05199_),
    .B2(\g_reduce0[4].adder.x[7] ),
    .ZN(_05235_));
 NAND3_X2 _28659_ (.A1(_05223_),
    .A2(_05167_),
    .A3(_05224_),
    .ZN(_05236_));
 NOR2_X1 _28660_ (.A1(_05116_),
    .A2(_05236_),
    .ZN(_05237_));
 AND2_X1 _28661_ (.A1(_05116_),
    .A2(_05236_),
    .ZN(_05238_));
 NOR2_X1 _28662_ (.A1(_05237_),
    .A2(_05238_),
    .ZN(_05239_));
 MUX2_X1 _28663_ (.A(_05230_),
    .B(_05239_),
    .S(_22262_),
    .Z(_05240_));
 OAI21_X1 _28664_ (.A(_05235_),
    .B1(_05240_),
    .B2(_05221_),
    .ZN(_00157_));
 OAI22_X2 _28665_ (.A1(\g_reduce0[6].adder.x[8] ),
    .A2(_05001_),
    .B1(_05208_),
    .B2(\g_reduce0[4].adder.x[8] ),
    .ZN(_05241_));
 NAND3_X1 _28666_ (.A1(_05228_),
    .A2(_05190_),
    .A3(_05193_),
    .ZN(_05242_));
 INV_X1 _28667_ (.A(_05116_),
    .ZN(_05243_));
 OR2_X1 _28668_ (.A1(_05243_),
    .A2(_05189_),
    .ZN(_05244_));
 XNOR2_X1 _28669_ (.A(_05091_),
    .B(_05244_),
    .ZN(_05245_));
 OR3_X1 _28670_ (.A1(_05228_),
    .A2(_05221_),
    .A3(_05245_),
    .ZN(_05246_));
 OAI211_X2 _28671_ (.A(_05238_),
    .B(_05242_),
    .C1(_05246_),
    .C2(_05190_),
    .ZN(_05247_));
 NAND2_X1 _28672_ (.A1(_05228_),
    .A2(_05193_),
    .ZN(_05248_));
 OAI21_X1 _28673_ (.A(_05246_),
    .B1(_05248_),
    .B2(_05237_),
    .ZN(_05249_));
 AOI21_X1 _28674_ (.A(_05241_),
    .B1(_05247_),
    .B2(_05249_),
    .ZN(_00158_));
 OAI22_X2 _28675_ (.A1(\g_reduce0[6].adder.x[9] ),
    .A2(_04585_),
    .B1(_05208_),
    .B2(\g_reduce0[4].adder.x[9] ),
    .ZN(_05250_));
 NAND2_X1 _28676_ (.A1(_05091_),
    .A2(_05116_),
    .ZN(_05251_));
 NOR4_X1 _28677_ (.A1(_05228_),
    .A2(_05251_),
    .A3(_05140_),
    .A4(_05236_),
    .ZN(_05252_));
 NAND3_X1 _28678_ (.A1(_05228_),
    .A2(_05091_),
    .A3(_05244_),
    .ZN(_05253_));
 NAND2_X1 _28679_ (.A1(_05251_),
    .A2(_05140_),
    .ZN(_05254_));
 OAI21_X1 _28680_ (.A(_05253_),
    .B1(_05254_),
    .B2(_05228_),
    .ZN(_05255_));
 NOR3_X1 _28681_ (.A1(_05221_),
    .A2(_05252_),
    .A3(_05255_),
    .ZN(_05256_));
 AND2_X1 _28682_ (.A1(_05167_),
    .A2(_05229_),
    .ZN(_05257_));
 NAND2_X1 _28683_ (.A1(_05140_),
    .A2(_05236_),
    .ZN(_05258_));
 NOR3_X1 _28684_ (.A1(_05228_),
    .A2(_05257_),
    .A3(_05258_),
    .ZN(_05259_));
 AOI21_X1 _28685_ (.A(_05244_),
    .B1(_05258_),
    .B2(_05091_),
    .ZN(_05260_));
 AOI21_X1 _28686_ (.A(_05259_),
    .B1(_05260_),
    .B2(_05228_),
    .ZN(_05261_));
 AOI21_X1 _28687_ (.A(_05250_),
    .B1(_05256_),
    .B2(_05261_),
    .ZN(_00159_));
 MUX2_X1 _28688_ (.A(_22265_),
    .B(\g_reduce0[4].adder.x[10] ),
    .S(_04589_),
    .Z(_05262_));
 MUX2_X1 _28689_ (.A(\g_reduce0[6].adder.x[10] ),
    .B(_05262_),
    .S(_05001_),
    .Z(_00145_));
 MUX2_X1 _28690_ (.A(_22273_),
    .B(_04581_),
    .S(_04589_),
    .Z(_05263_));
 MUX2_X1 _28691_ (.A(\g_reduce0[6].adder.x[11] ),
    .B(_05263_),
    .S(_05001_),
    .Z(_00146_));
 MUX2_X1 _28692_ (.A(_22138_),
    .B(_00584_),
    .S(_04629_),
    .Z(_05264_));
 NAND2_X1 _28693_ (.A1(_05017_),
    .A2(_22267_),
    .ZN(_05265_));
 XOR2_X1 _28694_ (.A(_05264_),
    .B(_05265_),
    .Z(_05266_));
 XNOR2_X1 _28695_ (.A(_14176_),
    .B(_22277_),
    .ZN(_05267_));
 MUX2_X1 _28696_ (.A(_05266_),
    .B(_05267_),
    .S(_05084_),
    .Z(_05268_));
 XOR2_X1 _28697_ (.A(_22272_),
    .B(_05268_),
    .Z(_05269_));
 MUX2_X1 _28698_ (.A(_04582_),
    .B(_05269_),
    .S(_05005_),
    .Z(_05270_));
 MUX2_X1 _28699_ (.A(\g_reduce0[6].adder.x[12] ),
    .B(_05270_),
    .S(_05001_),
    .Z(_00147_));
 MUX2_X1 _28700_ (.A(_22135_),
    .B(_00587_),
    .S(_04630_),
    .Z(_05271_));
 INV_X1 _28701_ (.A(_05271_),
    .ZN(_22278_));
 INV_X1 _28702_ (.A(_14173_),
    .ZN(_14178_));
 INV_X1 _28703_ (.A(_05264_),
    .ZN(_22274_));
 NAND4_X1 _28704_ (.A1(_05017_),
    .A2(_22266_),
    .A3(_14178_),
    .A4(_22274_),
    .ZN(_05272_));
 XNOR2_X1 _28705_ (.A(_22278_),
    .B(_05272_),
    .ZN(_05273_));
 INV_X1 _28706_ (.A(_22276_),
    .ZN(_05274_));
 INV_X1 _28707_ (.A(_14175_),
    .ZN(_05275_));
 AOI21_X1 _28708_ (.A(_22269_),
    .B1(_22270_),
    .B2(_05275_),
    .ZN(_05276_));
 INV_X1 _28709_ (.A(_22277_),
    .ZN(_05277_));
 OAI21_X1 _28710_ (.A(_05274_),
    .B1(_05276_),
    .B2(_05277_),
    .ZN(_05278_));
 XOR2_X1 _28711_ (.A(_22281_),
    .B(_05278_),
    .Z(_05279_));
 MUX2_X1 _28712_ (.A(_05273_),
    .B(_05279_),
    .S(_05084_),
    .Z(_05280_));
 NOR2_X1 _28713_ (.A1(_05017_),
    .A2(_14173_),
    .ZN(_05281_));
 AOI221_X2 _28714_ (.A(_05281_),
    .B1(_04981_),
    .B2(_05019_),
    .C1(_05017_),
    .C2(_22268_),
    .ZN(_05282_));
 AOI21_X2 _28715_ (.A(_05282_),
    .B1(_05084_),
    .B2(_14177_),
    .ZN(_22271_));
 NAND3_X1 _28716_ (.A1(_22264_),
    .A2(_05268_),
    .A3(_22271_),
    .ZN(_05283_));
 XNOR2_X1 _28717_ (.A(_05280_),
    .B(_05283_),
    .ZN(_05284_));
 MUX2_X1 _28718_ (.A(\g_reduce0[4].adder.x[13] ),
    .B(_05284_),
    .S(_05005_),
    .Z(_05285_));
 MUX2_X1 _28719_ (.A(\g_reduce0[6].adder.x[13] ),
    .B(_05285_),
    .S(_05001_),
    .Z(_00148_));
 NOR4_X1 _28720_ (.A1(_05084_),
    .A2(_05264_),
    .A3(_05265_),
    .A4(_05271_),
    .ZN(_05286_));
 OAI21_X1 _28721_ (.A(_05274_),
    .B1(_05277_),
    .B2(_14176_),
    .ZN(_05287_));
 AOI21_X1 _28722_ (.A(_22280_),
    .B1(_05287_),
    .B2(_22281_),
    .ZN(_05288_));
 AOI21_X1 _28723_ (.A(_05286_),
    .B1(_05288_),
    .B2(_05084_),
    .ZN(_05289_));
 NAND3_X1 _28724_ (.A1(_22272_),
    .A2(_05268_),
    .A3(_05280_),
    .ZN(_05290_));
 XOR2_X1 _28725_ (.A(_05289_),
    .B(_05290_),
    .Z(_05291_));
 AND3_X1 _28726_ (.A1(_04586_),
    .A2(_04603_),
    .A3(_05291_),
    .ZN(_05292_));
 OAI21_X1 _28727_ (.A(_05005_),
    .B1(_04603_),
    .B2(_05291_),
    .ZN(_05293_));
 OAI21_X1 _28728_ (.A(_04583_),
    .B1(_05292_),
    .B2(_05293_),
    .ZN(_05294_));
 NAND2_X1 _28729_ (.A1(\g_reduce0[6].adder.x[14] ),
    .A2(_04603_),
    .ZN(_05295_));
 NOR2_X1 _28730_ (.A1(_05291_),
    .A2(_05295_),
    .ZN(_05296_));
 OAI21_X1 _28731_ (.A(_05295_),
    .B1(_04585_),
    .B2(\g_reduce0[6].adder.x[14] ),
    .ZN(_05297_));
 NOR2_X1 _28732_ (.A1(_04583_),
    .A2(_05297_),
    .ZN(_05298_));
 AOI21_X1 _28733_ (.A(_05296_),
    .B1(_05298_),
    .B2(_05291_),
    .ZN(_05299_));
 OAI221_X2 _28734_ (.A(_05294_),
    .B1(_05299_),
    .B2(_04589_),
    .C1(_05001_),
    .C2(_04586_),
    .ZN(_00149_));
 BUF_X2 _28735_ (.A(\g_reduce0[8].adder.x[11] ),
    .Z(_05300_));
 BUF_X2 _28736_ (.A(\g_reduce0[8].adder.x[12] ),
    .Z(_05301_));
 BUF_X2 _28737_ (.A(\g_reduce0[8].adder.x[14] ),
    .Z(_05302_));
 OR2_X1 _28738_ (.A1(\g_reduce0[8].adder.x[10] ),
    .A2(\g_reduce0[8].adder.x[13] ),
    .ZN(_05303_));
 NOR4_X4 _28739_ (.A1(_05300_),
    .A2(_05301_),
    .A3(_05302_),
    .A4(_05303_),
    .ZN(_05304_));
 BUF_X2 _28740_ (.A(\g_reduce0[10].adder.x[14] ),
    .Z(_05305_));
 OR2_X1 _28741_ (.A1(\g_reduce0[10].adder.x[10] ),
    .A2(\g_reduce0[10].adder.x[13] ),
    .ZN(_05306_));
 OR4_X2 _28742_ (.A1(\g_reduce0[10].adder.x[11] ),
    .A2(\g_reduce0[10].adder.x[12] ),
    .A3(_05305_),
    .A4(_05306_),
    .ZN(_05307_));
 CLKBUF_X3 _28743_ (.A(_05307_),
    .Z(_05308_));
 INV_X1 _28744_ (.A(_22328_),
    .ZN(_05309_));
 INV_X1 _28745_ (.A(_22286_),
    .ZN(_05310_));
 INV_X1 _28746_ (.A(_22322_),
    .ZN(_05311_));
 AOI21_X1 _28747_ (.A(_22289_),
    .B1(_05311_),
    .B2(_22290_),
    .ZN(_05312_));
 BUF_X2 _28748_ (.A(_22287_),
    .Z(_05313_));
 INV_X1 _28749_ (.A(_05313_),
    .ZN(_05314_));
 OAI21_X1 _28750_ (.A(_05310_),
    .B1(_05312_),
    .B2(_05314_),
    .ZN(_05315_));
 BUF_X4 _28751_ (.A(_22284_),
    .Z(_05316_));
 AOI21_X2 _28752_ (.A(_22283_),
    .B1(_05315_),
    .B2(_05316_),
    .ZN(_05317_));
 INV_X4 _28753_ (.A(_22329_),
    .ZN(_05318_));
 OAI21_X4 _28754_ (.A(_05309_),
    .B1(_05317_),
    .B2(_05318_),
    .ZN(_05319_));
 BUF_X2 _28755_ (.A(_22323_),
    .Z(_05320_));
 INV_X2 _28756_ (.A(_05320_),
    .ZN(_05321_));
 INV_X1 _28757_ (.A(_22290_),
    .ZN(_05322_));
 NAND2_X2 _28758_ (.A1(_05316_),
    .A2(_05313_),
    .ZN(_05323_));
 OR4_X1 _28759_ (.A1(_05318_),
    .A2(_05321_),
    .A3(_05322_),
    .A4(_05323_),
    .ZN(_05324_));
 BUF_X4 _28760_ (.A(_05324_),
    .Z(_05325_));
 INV_X1 _28761_ (.A(_22295_),
    .ZN(_05326_));
 AOI21_X1 _28762_ (.A(_22298_),
    .B1(_22299_),
    .B2(_22301_),
    .ZN(_05327_));
 INV_X1 _28763_ (.A(_22296_),
    .ZN(_05328_));
 OAI21_X2 _28764_ (.A(_05326_),
    .B1(_05327_),
    .B2(_05328_),
    .ZN(_05329_));
 AOI21_X2 _28765_ (.A(_22292_),
    .B1(_05329_),
    .B2(_22293_),
    .ZN(_05330_));
 NAND3_X2 _28766_ (.A1(_22305_),
    .A2(_22308_),
    .A3(_22311_),
    .ZN(_05331_));
 INV_X1 _28767_ (.A(_05331_),
    .ZN(_05332_));
 INV_X1 _28768_ (.A(_22313_),
    .ZN(_05333_));
 INV_X1 _28769_ (.A(_22314_),
    .ZN(_05334_));
 INV_X1 _28770_ (.A(_22319_),
    .ZN(_05335_));
 AOI21_X1 _28771_ (.A(_22316_),
    .B1(_05335_),
    .B2(_22317_),
    .ZN(_05336_));
 OAI21_X1 _28772_ (.A(_05333_),
    .B1(_05334_),
    .B2(_05336_),
    .ZN(_05337_));
 AND2_X1 _28773_ (.A1(_22308_),
    .A2(_22310_),
    .ZN(_05338_));
 OR2_X1 _28774_ (.A1(_22307_),
    .A2(_05338_),
    .ZN(_05339_));
 AOI221_X2 _28775_ (.A(_22304_),
    .B1(_05332_),
    .B2(_05337_),
    .C1(_05339_),
    .C2(_22305_),
    .ZN(_05340_));
 NAND4_X4 _28776_ (.A1(_22293_),
    .A2(_22296_),
    .A3(_22299_),
    .A4(_22302_),
    .ZN(_05341_));
 OAI21_X4 _28777_ (.A(_05330_),
    .B1(_05340_),
    .B2(_05341_),
    .ZN(_05342_));
 NAND3_X2 _28778_ (.A1(_22314_),
    .A2(_22317_),
    .A3(_22320_),
    .ZN(_05343_));
 NOR3_X4 _28779_ (.A1(_05341_),
    .A2(_05331_),
    .A3(_05343_),
    .ZN(_05344_));
 NOR2_X1 _28780_ (.A1(_05325_),
    .A2(_05344_),
    .ZN(_05345_));
 AOI22_X4 _28781_ (.A1(_05319_),
    .A2(_05325_),
    .B1(_05342_),
    .B2(_05345_),
    .ZN(_05346_));
 AOI21_X1 _28782_ (.A(_05304_),
    .B1(_05308_),
    .B2(_05346_),
    .ZN(_05347_));
 MUX2_X1 _28783_ (.A(\g_reduce0[10].adder.x[15] ),
    .B(\g_reduce0[8].adder.x[15] ),
    .S(_05347_),
    .Z(_00166_));
 INV_X1 _28784_ (.A(_22283_),
    .ZN(_05348_));
 INV_X1 _28785_ (.A(_22289_),
    .ZN(_05349_));
 OAI21_X1 _28786_ (.A(_05349_),
    .B1(_22322_),
    .B2(_05322_),
    .ZN(_05350_));
 AOI21_X1 _28787_ (.A(_22286_),
    .B1(_05350_),
    .B2(_05313_),
    .ZN(_05351_));
 INV_X2 _28788_ (.A(_05316_),
    .ZN(_05352_));
 OAI21_X2 _28789_ (.A(_05348_),
    .B1(_05351_),
    .B2(_05352_),
    .ZN(_05353_));
 AOI21_X4 _28790_ (.A(_22328_),
    .B1(_05353_),
    .B2(_22329_),
    .ZN(_05354_));
 NOR4_X4 _28791_ (.A1(_05318_),
    .A2(_05321_),
    .A3(_05322_),
    .A4(_05323_),
    .ZN(_05355_));
 INV_X1 _28792_ (.A(_05341_),
    .ZN(_05356_));
 AOI21_X1 _28793_ (.A(_22304_),
    .B1(_05339_),
    .B2(_22305_),
    .ZN(_05357_));
 INV_X1 _28794_ (.A(_22316_),
    .ZN(_05358_));
 INV_X1 _28795_ (.A(_22317_),
    .ZN(_05359_));
 OAI21_X1 _28796_ (.A(_05358_),
    .B1(_22319_),
    .B2(_05359_),
    .ZN(_05360_));
 AOI21_X1 _28797_ (.A(_22313_),
    .B1(_22314_),
    .B2(_05360_),
    .ZN(_05361_));
 OAI21_X1 _28798_ (.A(_05357_),
    .B1(_05361_),
    .B2(_05331_),
    .ZN(_05362_));
 AOI221_X2 _28799_ (.A(_22292_),
    .B1(_05356_),
    .B2(_05362_),
    .C1(_05329_),
    .C2(_22293_),
    .ZN(_05363_));
 OR2_X2 _28800_ (.A1(_05325_),
    .A2(_05344_),
    .ZN(_05364_));
 OAI22_X4 _28801_ (.A1(_05354_),
    .A2(_05355_),
    .B1(_05363_),
    .B2(_05364_),
    .ZN(_05365_));
 BUF_X8 _28802_ (.A(_05365_),
    .Z(_05366_));
 BUF_X8 _28803_ (.A(_05366_),
    .Z(_05367_));
 MUX2_X2 _28804_ (.A(_00590_),
    .B(_22321_),
    .S(_05367_),
    .Z(_22407_));
 NOR2_X2 _28805_ (.A1(_05301_),
    .A2(_22285_),
    .ZN(_05368_));
 NOR2_X1 _28806_ (.A1(_05300_),
    .A2(_22288_),
    .ZN(_05369_));
 BUF_X2 _28807_ (.A(_05313_),
    .Z(_05370_));
 AOI21_X1 _28808_ (.A(_05368_),
    .B1(_05369_),
    .B2(_05370_),
    .ZN(_05371_));
 NOR2_X2 _28809_ (.A1(\g_reduce0[10].adder.x[12] ),
    .A2(_00598_),
    .ZN(_05372_));
 NOR2_X1 _28810_ (.A1(\g_reduce0[10].adder.x[11] ),
    .A2(_00593_),
    .ZN(_05373_));
 AOI21_X1 _28811_ (.A(_05372_),
    .B1(_05373_),
    .B2(_05370_),
    .ZN(_05374_));
 MUX2_X2 _28812_ (.A(_05371_),
    .B(_05374_),
    .S(_05366_),
    .Z(_05375_));
 NAND2_X1 _28813_ (.A1(_05370_),
    .A2(_22290_),
    .ZN(_05376_));
 INV_X1 _28814_ (.A(_22321_),
    .ZN(_05377_));
 NOR2_X2 _28815_ (.A1(_00590_),
    .A2(_05377_),
    .ZN(_05378_));
 AND3_X1 _28816_ (.A1(_05342_),
    .A2(_05345_),
    .A3(_05378_),
    .ZN(_05379_));
 AND3_X1 _28817_ (.A1(_05319_),
    .A2(_05325_),
    .A3(_05378_),
    .ZN(_05380_));
 NAND2_X1 _28818_ (.A1(_00590_),
    .A2(_05377_),
    .ZN(_05381_));
 AOI221_X2 _28819_ (.A(_05381_),
    .B1(_05345_),
    .B2(_05342_),
    .C1(_05319_),
    .C2(_05325_),
    .ZN(_05382_));
 OR4_X4 _28820_ (.A1(_05376_),
    .A2(_05379_),
    .A3(_05380_),
    .A4(_05382_),
    .ZN(_05383_));
 AOI21_X4 _28821_ (.A(_05352_),
    .B1(_05375_),
    .B2(_05383_),
    .ZN(_05384_));
 INV_X1 _28822_ (.A(_05371_),
    .ZN(_05385_));
 INV_X1 _28823_ (.A(_05374_),
    .ZN(_05386_));
 MUX2_X2 _28824_ (.A(_05385_),
    .B(_05386_),
    .S(_05365_),
    .Z(_05387_));
 AOI211_X2 _28825_ (.A(_05376_),
    .B(_05382_),
    .C1(_05378_),
    .C2(_05365_),
    .ZN(_05388_));
 NOR3_X4 _28826_ (.A1(_05316_),
    .A2(_05387_),
    .A3(_05388_),
    .ZN(_05389_));
 NOR2_X4 _28827_ (.A1(_05384_),
    .A2(_05389_),
    .ZN(_05390_));
 NOR2_X1 _28828_ (.A1(\g_reduce0[10].adder.x[13] ),
    .A2(_00601_),
    .ZN(_05391_));
 AOI21_X1 _28829_ (.A(_05391_),
    .B1(_05372_),
    .B2(_05316_),
    .ZN(_05392_));
 OR2_X1 _28830_ (.A1(_05346_),
    .A2(_05392_),
    .ZN(_05393_));
 NOR2_X1 _28831_ (.A1(_22325_),
    .A2(_05369_),
    .ZN(_05394_));
 NOR2_X1 _28832_ (.A1(_22325_),
    .A2(_05373_),
    .ZN(_05395_));
 MUX2_X1 _28833_ (.A(_05394_),
    .B(_05395_),
    .S(_05366_),
    .Z(_05396_));
 NOR2_X1 _28834_ (.A1(\g_reduce0[8].adder.x[13] ),
    .A2(_22282_),
    .ZN(_05397_));
 AOI21_X1 _28835_ (.A(_05397_),
    .B1(_05368_),
    .B2(_05316_),
    .ZN(_05398_));
 OAI221_X2 _28836_ (.A(_05393_),
    .B1(_05396_),
    .B2(_05323_),
    .C1(_05367_),
    .C2(_05398_),
    .ZN(_05399_));
 XNOR2_X2 _28837_ (.A(_05318_),
    .B(_05399_),
    .ZN(_05400_));
 OR2_X1 _28838_ (.A1(_05390_),
    .A2(_05400_),
    .ZN(_05401_));
 MUX2_X1 _28839_ (.A(_00596_),
    .B(_22297_),
    .S(_05367_),
    .Z(_05402_));
 MUX2_X1 _28840_ (.A(_00597_),
    .B(_22300_),
    .S(_05367_),
    .Z(_05403_));
 CLKBUF_X3 _28841_ (.A(_05320_),
    .Z(_05404_));
 MUX2_X1 _28842_ (.A(_05402_),
    .B(_05403_),
    .S(_05404_),
    .Z(_05405_));
 CLKBUF_X3 _28843_ (.A(_05367_),
    .Z(_05406_));
 MUX2_X1 _28844_ (.A(_00594_),
    .B(_22303_),
    .S(_05406_),
    .Z(_05407_));
 MUX2_X1 _28845_ (.A(_00595_),
    .B(_22306_),
    .S(_05406_),
    .Z(_05408_));
 MUX2_X1 _28846_ (.A(_05407_),
    .B(_05408_),
    .S(_05404_),
    .Z(_05409_));
 CLKBUF_X3 _28847_ (.A(_22326_),
    .Z(_05410_));
 INV_X2 _28848_ (.A(_05410_),
    .ZN(_05411_));
 MUX2_X1 _28849_ (.A(_05405_),
    .B(_05409_),
    .S(_05411_),
    .Z(_05412_));
 MUX2_X1 _28850_ (.A(_00591_),
    .B(_22309_),
    .S(_05406_),
    .Z(_05413_));
 MUX2_X1 _28851_ (.A(_00592_),
    .B(_22312_),
    .S(_05406_),
    .Z(_05414_));
 MUX2_X1 _28852_ (.A(_05413_),
    .B(_05414_),
    .S(_05404_),
    .Z(_05415_));
 MUX2_X1 _28853_ (.A(_22318_),
    .B(_00589_),
    .S(_05366_),
    .Z(_05416_));
 MUX2_X1 _28854_ (.A(_00588_),
    .B(_22315_),
    .S(_05406_),
    .Z(_05417_));
 MUX2_X1 _28855_ (.A(_05416_),
    .B(_05417_),
    .S(_05321_),
    .Z(_05418_));
 MUX2_X1 _28856_ (.A(_05415_),
    .B(_05418_),
    .S(_05411_),
    .Z(_05419_));
 NOR2_X1 _28857_ (.A1(_05314_),
    .A2(_05395_),
    .ZN(_05420_));
 OR2_X1 _28858_ (.A1(_22325_),
    .A2(_05373_),
    .ZN(_05421_));
 NOR2_X1 _28859_ (.A1(_05370_),
    .A2(_05421_),
    .ZN(_05422_));
 OAI21_X2 _28860_ (.A(_05366_),
    .B1(_05420_),
    .B2(_05422_),
    .ZN(_05423_));
 NOR2_X1 _28861_ (.A1(_05314_),
    .A2(_05394_),
    .ZN(_05424_));
 OR2_X1 _28862_ (.A1(_22325_),
    .A2(_05369_),
    .ZN(_05425_));
 NOR2_X1 _28863_ (.A1(_05370_),
    .A2(_05425_),
    .ZN(_05426_));
 OAI21_X2 _28864_ (.A(_05346_),
    .B1(_05424_),
    .B2(_05426_),
    .ZN(_05427_));
 NAND2_X2 _28865_ (.A1(_05423_),
    .A2(_05427_),
    .ZN(_05428_));
 MUX2_X1 _28866_ (.A(_05412_),
    .B(_05419_),
    .S(_05428_),
    .Z(_05429_));
 MUX2_X1 _28867_ (.A(_00600_),
    .B(_22294_),
    .S(_05367_),
    .Z(_05430_));
 OR2_X1 _28868_ (.A1(_05321_),
    .A2(_05430_),
    .ZN(_05431_));
 MUX2_X1 _28869_ (.A(_00599_),
    .B(_22291_),
    .S(_05406_),
    .Z(_05432_));
 OAI21_X1 _28870_ (.A(_05431_),
    .B1(_05432_),
    .B2(_05404_),
    .ZN(_05433_));
 MUX2_X1 _28871_ (.A(_05404_),
    .B(_05433_),
    .S(_05411_),
    .Z(_05434_));
 NAND2_X1 _28872_ (.A1(_05428_),
    .A2(_05434_),
    .ZN(_05435_));
 NOR2_X1 _28873_ (.A1(_05370_),
    .A2(_05368_),
    .ZN(_05436_));
 OAI221_X2 _28874_ (.A(_05436_),
    .B1(_05364_),
    .B2(_05363_),
    .C1(_05354_),
    .C2(_05355_),
    .ZN(_05437_));
 OR2_X1 _28875_ (.A1(_05370_),
    .A2(_05372_),
    .ZN(_05438_));
 OAI211_X2 _28876_ (.A(_05316_),
    .B(_05437_),
    .C1(_05438_),
    .C2(_05346_),
    .ZN(_05439_));
 INV_X1 _28877_ (.A(_05397_),
    .ZN(_05440_));
 INV_X1 _28878_ (.A(_05391_),
    .ZN(_05441_));
 MUX2_X1 _28879_ (.A(_05440_),
    .B(_05441_),
    .S(_05366_),
    .Z(_05442_));
 AOI21_X2 _28880_ (.A(_05318_),
    .B1(_05439_),
    .B2(_05442_),
    .ZN(_05443_));
 OR2_X1 _28881_ (.A1(_05313_),
    .A2(_05368_),
    .ZN(_05444_));
 AOI221_X2 _28882_ (.A(_05444_),
    .B1(_05345_),
    .B2(_05342_),
    .C1(_05319_),
    .C2(_05325_),
    .ZN(_05445_));
 NOR2_X1 _28883_ (.A1(_05370_),
    .A2(_05372_),
    .ZN(_05446_));
 AOI211_X2 _28884_ (.A(_05352_),
    .B(_05445_),
    .C1(_05446_),
    .C2(_05365_),
    .ZN(_05447_));
 MUX2_X2 _28885_ (.A(_05397_),
    .B(_05391_),
    .S(_05365_),
    .Z(_05448_));
 NOR3_X4 _28886_ (.A1(_22329_),
    .A2(_05447_),
    .A3(_05448_),
    .ZN(_05449_));
 OAI21_X1 _28887_ (.A(_05390_),
    .B1(_05443_),
    .B2(_05449_),
    .ZN(_05450_));
 OAI22_X2 _28888_ (.A1(_05401_),
    .A2(_05429_),
    .B1(_05435_),
    .B2(_05450_),
    .ZN(_22390_));
 AOI21_X1 _28889_ (.A(_05410_),
    .B1(_05432_),
    .B2(_05404_),
    .ZN(_05451_));
 NAND2_X1 _28890_ (.A1(_05428_),
    .A2(_05451_),
    .ZN(_05452_));
 MUX2_X1 _28891_ (.A(_00597_),
    .B(_00594_),
    .S(_05320_),
    .Z(_05453_));
 AOI221_X2 _28892_ (.A(_05453_),
    .B1(_05345_),
    .B2(_05342_),
    .C1(_05319_),
    .C2(_05325_),
    .ZN(_05454_));
 MUX2_X1 _28893_ (.A(_22300_),
    .B(_22303_),
    .S(_05320_),
    .Z(_05455_));
 INV_X1 _28894_ (.A(_05455_),
    .ZN(_05456_));
 AOI21_X1 _28895_ (.A(_05454_),
    .B1(_05456_),
    .B2(_05406_),
    .ZN(_05457_));
 MUX2_X1 _28896_ (.A(_05402_),
    .B(_05430_),
    .S(_05321_),
    .Z(_05458_));
 MUX2_X1 _28897_ (.A(_05457_),
    .B(_05458_),
    .S(_05410_),
    .Z(_05459_));
 MUX2_X1 _28898_ (.A(_00595_),
    .B(_00591_),
    .S(_05320_),
    .Z(_05460_));
 AOI221_X2 _28899_ (.A(_05460_),
    .B1(_05345_),
    .B2(_05342_),
    .C1(_05319_),
    .C2(_05325_),
    .ZN(_05461_));
 MUX2_X1 _28900_ (.A(_22306_),
    .B(_22309_),
    .S(_05320_),
    .Z(_05462_));
 INV_X1 _28901_ (.A(_05462_),
    .ZN(_05463_));
 AOI21_X1 _28902_ (.A(_05461_),
    .B1(_05463_),
    .B2(_05406_),
    .ZN(_05464_));
 MUX2_X1 _28903_ (.A(_00592_),
    .B(_00588_),
    .S(_05320_),
    .Z(_05465_));
 MUX2_X1 _28904_ (.A(_22312_),
    .B(_22315_),
    .S(_05404_),
    .Z(_05466_));
 MUX2_X1 _28905_ (.A(_05465_),
    .B(_05466_),
    .S(_05366_),
    .Z(_05467_));
 MUX2_X1 _28906_ (.A(_05464_),
    .B(_05467_),
    .S(_05411_),
    .Z(_05468_));
 MUX2_X1 _28907_ (.A(_05459_),
    .B(_05468_),
    .S(_05428_),
    .Z(_05469_));
 OAI21_X4 _28908_ (.A(_05316_),
    .B1(_05387_),
    .B2(_05388_),
    .ZN(_05470_));
 NAND3_X4 _28909_ (.A1(_05352_),
    .A2(_05375_),
    .A3(_05383_),
    .ZN(_05471_));
 NAND2_X2 _28910_ (.A1(_05470_),
    .A2(_05471_),
    .ZN(_05472_));
 MUX2_X1 _28911_ (.A(_05452_),
    .B(_05469_),
    .S(_05472_),
    .Z(_05473_));
 OR2_X1 _28912_ (.A1(_05400_),
    .A2(_05473_),
    .ZN(_14186_));
 INV_X1 _28913_ (.A(_14186_),
    .ZN(_14180_));
 INV_X1 _28914_ (.A(_22390_),
    .ZN(_22393_));
 OR2_X1 _28915_ (.A1(_05401_),
    .A2(_05452_),
    .ZN(_22345_));
 INV_X1 _28916_ (.A(_22345_),
    .ZN(_22349_));
 NOR2_X2 _28917_ (.A1(_05390_),
    .A2(_05400_),
    .ZN(_05474_));
 NAND3_X1 _28918_ (.A1(_05474_),
    .A2(_05428_),
    .A3(_05434_),
    .ZN(_22339_));
 INV_X1 _28919_ (.A(_22339_),
    .ZN(_22342_));
 MUX2_X1 _28920_ (.A(_00596_),
    .B(_00599_),
    .S(_05410_),
    .Z(_05475_));
 NOR2_X1 _28921_ (.A1(_05404_),
    .A2(_05410_),
    .ZN(_05476_));
 AOI22_X1 _28922_ (.A1(_05404_),
    .A2(_05475_),
    .B1(_05476_),
    .B2(_00600_),
    .ZN(_05477_));
 MUX2_X1 _28923_ (.A(_22297_),
    .B(_22291_),
    .S(_05410_),
    .Z(_05478_));
 AOI22_X1 _28924_ (.A1(_22294_),
    .A2(_05476_),
    .B1(_05478_),
    .B2(_05404_),
    .ZN(_05479_));
 MUX2_X1 _28925_ (.A(_05477_),
    .B(_05479_),
    .S(_05367_),
    .Z(_05480_));
 NAND2_X1 _28926_ (.A1(_05370_),
    .A2(_05425_),
    .ZN(_05481_));
 NAND2_X1 _28927_ (.A1(_05314_),
    .A2(_05394_),
    .ZN(_05482_));
 AOI21_X4 _28928_ (.A(_05366_),
    .B1(_05481_),
    .B2(_05482_),
    .ZN(_05483_));
 NAND2_X1 _28929_ (.A1(_05370_),
    .A2(_05421_),
    .ZN(_05484_));
 NAND2_X1 _28930_ (.A1(_05314_),
    .A2(_05395_),
    .ZN(_05485_));
 AOI21_X4 _28931_ (.A(_05346_),
    .B1(_05484_),
    .B2(_05485_),
    .ZN(_05486_));
 OAI21_X1 _28932_ (.A(_05480_),
    .B1(_05483_),
    .B2(_05486_),
    .ZN(_05487_));
 OR2_X1 _28933_ (.A1(_05401_),
    .A2(_05487_),
    .ZN(_22373_));
 INV_X1 _28934_ (.A(_22373_),
    .ZN(_22377_));
 NOR2_X1 _28935_ (.A1(_05411_),
    .A2(_05433_),
    .ZN(_05488_));
 AOI21_X1 _28936_ (.A(_05488_),
    .B1(_05405_),
    .B2(_05411_),
    .ZN(_05489_));
 NOR2_X2 _28937_ (.A1(_05321_),
    .A2(_05410_),
    .ZN(_05490_));
 NOR2_X4 _28938_ (.A1(_05486_),
    .A2(_05483_),
    .ZN(_05491_));
 MUX2_X1 _28939_ (.A(_05489_),
    .B(_05490_),
    .S(_05491_),
    .Z(_05492_));
 NAND2_X1 _28940_ (.A1(_05474_),
    .A2(_05492_),
    .ZN(_22353_));
 INV_X1 _28941_ (.A(_22353_),
    .ZN(_22356_));
 NOR2_X1 _28942_ (.A1(_05491_),
    .A2(_05459_),
    .ZN(_05493_));
 AOI21_X1 _28943_ (.A(_05493_),
    .B1(_05451_),
    .B2(_05491_),
    .ZN(_05494_));
 NOR2_X1 _28944_ (.A1(_05401_),
    .A2(_05494_),
    .ZN(_22360_));
 INV_X1 _28945_ (.A(_22360_),
    .ZN(_22363_));
 NAND2_X1 _28946_ (.A1(_05491_),
    .A2(_05434_),
    .ZN(_05495_));
 OAI21_X1 _28947_ (.A(_05495_),
    .B1(_05491_),
    .B2(_05412_),
    .ZN(_05496_));
 AND2_X1 _28948_ (.A1(_05474_),
    .A2(_05496_),
    .ZN(_22366_));
 INV_X1 _28949_ (.A(_22366_),
    .ZN(_22370_));
 NAND2_X1 _28950_ (.A1(_05491_),
    .A2(_05480_),
    .ZN(_05497_));
 AOI211_X2 _28951_ (.A(_05411_),
    .B(_05454_),
    .C1(_05456_),
    .C2(_05366_),
    .ZN(_05498_));
 AOI211_X2 _28952_ (.A(_05410_),
    .B(_05461_),
    .C1(_05463_),
    .C2(_05366_),
    .ZN(_05499_));
 OR2_X1 _28953_ (.A1(_05498_),
    .A2(_05499_),
    .ZN(_05500_));
 OAI21_X1 _28954_ (.A(_05497_),
    .B1(_05500_),
    .B2(_05491_),
    .ZN(_05501_));
 AND2_X1 _28955_ (.A1(_05474_),
    .A2(_05501_),
    .ZN(_22383_));
 INV_X1 _28956_ (.A(_22383_),
    .ZN(_22387_));
 OAI21_X2 _28957_ (.A(_05490_),
    .B1(_05483_),
    .B2(_05486_),
    .ZN(_05502_));
 NAND3_X2 _28958_ (.A1(_05318_),
    .A2(_05439_),
    .A3(_05442_),
    .ZN(_05503_));
 OAI21_X2 _28959_ (.A(_22329_),
    .B1(_05447_),
    .B2(_05448_),
    .ZN(_05504_));
 AOI21_X4 _28960_ (.A(_05502_),
    .B1(_05503_),
    .B2(_05504_),
    .ZN(_05505_));
 NAND2_X1 _28961_ (.A1(_05491_),
    .A2(_05489_),
    .ZN(_05506_));
 MUX2_X1 _28962_ (.A(_05409_),
    .B(_05415_),
    .S(_05411_),
    .Z(_05507_));
 OAI21_X1 _28963_ (.A(_05506_),
    .B1(_05507_),
    .B2(_05491_),
    .ZN(_05508_));
 AOI22_X2 _28964_ (.A1(_05390_),
    .A2(_05505_),
    .B1(_05508_),
    .B2(_05474_),
    .ZN(_22380_));
 INV_X1 _28965_ (.A(_22380_),
    .ZN(_22334_));
 XNOR2_X2 _28966_ (.A(\g_reduce0[10].adder.x[15] ),
    .B(\g_reduce0[8].adder.x[15] ),
    .ZN(_05509_));
 CLKBUF_X3 _28967_ (.A(_05509_),
    .Z(_05510_));
 CLKBUF_X3 _28968_ (.A(_22348_),
    .Z(_05511_));
 BUF_X2 _28969_ (.A(_22341_),
    .Z(_05512_));
 OR2_X1 _28970_ (.A1(_22378_),
    .A2(_22357_),
    .ZN(_05513_));
 OR3_X1 _28971_ (.A1(_22361_),
    .A2(_22368_),
    .A3(_05513_),
    .ZN(_05514_));
 INV_X1 _28972_ (.A(_22385_),
    .ZN(_05515_));
 BUF_X1 _28973_ (.A(_22337_),
    .Z(_05516_));
 AOI21_X1 _28974_ (.A(_22336_),
    .B1(_14183_),
    .B2(_05516_),
    .ZN(_05517_));
 BUF_X2 _28975_ (.A(_22386_),
    .Z(_05518_));
 INV_X1 _28976_ (.A(_05518_),
    .ZN(_05519_));
 OAI21_X2 _28977_ (.A(_05515_),
    .B1(_05517_),
    .B2(_05519_),
    .ZN(_05520_));
 CLKBUF_X3 _28978_ (.A(_22369_),
    .Z(_05521_));
 AOI21_X2 _28979_ (.A(_05514_),
    .B1(_05520_),
    .B2(_05521_),
    .ZN(_05522_));
 INV_X1 _28980_ (.A(_22378_),
    .ZN(_05523_));
 BUF_X2 _28981_ (.A(_22376_),
    .Z(_05524_));
 NAND2_X1 _28982_ (.A1(_05523_),
    .A2(_05524_),
    .ZN(_05525_));
 CLKBUF_X2 _28983_ (.A(_22355_),
    .Z(_05526_));
 BUF_X2 _28984_ (.A(_22362_),
    .Z(_05527_));
 INV_X2 _28985_ (.A(_05527_),
    .ZN(_05528_));
 INV_X1 _28986_ (.A(_22361_),
    .ZN(_05529_));
 AOI21_X2 _28987_ (.A(_05526_),
    .B1(_05528_),
    .B2(_05529_),
    .ZN(_05530_));
 OAI21_X1 _28988_ (.A(_05525_),
    .B1(_05513_),
    .B2(_05530_),
    .ZN(_05531_));
 OR3_X1 _28989_ (.A1(_05512_),
    .A2(_05522_),
    .A3(_05531_),
    .ZN(_05532_));
 INV_X1 _28990_ (.A(_22343_),
    .ZN(_05533_));
 AOI21_X1 _28991_ (.A(_05511_),
    .B1(_05532_),
    .B2(_05533_),
    .ZN(_05534_));
 OAI21_X2 _28992_ (.A(_05510_),
    .B1(_05534_),
    .B2(_22350_),
    .ZN(_05535_));
 INV_X1 _28993_ (.A(_05511_),
    .ZN(_05536_));
 INV_X1 _28994_ (.A(_22340_),
    .ZN(_05537_));
 INV_X1 _28995_ (.A(_22375_),
    .ZN(_05538_));
 OAI21_X1 _28996_ (.A(_05524_),
    .B1(_22354_),
    .B2(_05526_),
    .ZN(_05539_));
 NAND2_X1 _28997_ (.A1(_05538_),
    .A2(_05539_),
    .ZN(_05540_));
 AOI21_X2 _28998_ (.A(_22381_),
    .B1(_14187_),
    .B2(_22382_),
    .ZN(_05541_));
 OR4_X2 _28999_ (.A1(_05527_),
    .A2(_05521_),
    .A3(_05518_),
    .A4(_05541_),
    .ZN(_05542_));
 NOR2_X1 _29000_ (.A1(_05527_),
    .A2(_05521_),
    .ZN(_05543_));
 AOI221_X2 _29001_ (.A(_22364_),
    .B1(_05528_),
    .B2(_22371_),
    .C1(_22388_),
    .C2(_05543_),
    .ZN(_05544_));
 NOR2_X1 _29002_ (.A1(_22375_),
    .A2(_22354_),
    .ZN(_05545_));
 NAND3_X1 _29003_ (.A1(_05542_),
    .A2(_05544_),
    .A3(_05545_),
    .ZN(_05546_));
 NAND3_X1 _29004_ (.A1(_05512_),
    .A2(_05540_),
    .A3(_05546_),
    .ZN(_05547_));
 AOI21_X1 _29005_ (.A(_05536_),
    .B1(_05537_),
    .B2(_05547_),
    .ZN(_05548_));
 OR3_X2 _29006_ (.A1(_22347_),
    .A2(_05510_),
    .A3(_05548_),
    .ZN(_05549_));
 NAND2_X4 _29007_ (.A1(_05535_),
    .A2(_05549_),
    .ZN(_05550_));
 NOR2_X1 _29008_ (.A1(_05523_),
    .A2(_05512_),
    .ZN(_05551_));
 OAI21_X1 _29009_ (.A(_05509_),
    .B1(_05551_),
    .B2(_22343_),
    .ZN(_05552_));
 XOR2_X2 _29010_ (.A(\g_reduce0[10].adder.x[15] ),
    .B(\g_reduce0[8].adder.x[15] ),
    .Z(_05553_));
 OR3_X1 _29011_ (.A1(_05512_),
    .A2(_05524_),
    .A3(_05553_),
    .ZN(_05554_));
 NOR2_X1 _29012_ (.A1(_22361_),
    .A2(_22368_),
    .ZN(_05555_));
 AOI21_X2 _29013_ (.A(_22330_),
    .B1(_14181_),
    .B2(_22331_),
    .ZN(_05556_));
 NAND3_X1 _29014_ (.A1(_05521_),
    .A2(_05518_),
    .A3(_05516_),
    .ZN(_05557_));
 AOI21_X2 _29015_ (.A(_22385_),
    .B1(_05518_),
    .B2(_22336_),
    .ZN(_05558_));
 INV_X1 _29016_ (.A(_05521_),
    .ZN(_05559_));
 OAI221_X2 _29017_ (.A(_05555_),
    .B1(_05556_),
    .B2(_05557_),
    .C1(_05558_),
    .C2(_05559_),
    .ZN(_05560_));
 AOI21_X2 _29018_ (.A(_22357_),
    .B1(_05530_),
    .B2(_05560_),
    .ZN(_05561_));
 OAI21_X1 _29019_ (.A(_05552_),
    .B1(_05554_),
    .B2(_05561_),
    .ZN(_05562_));
 NAND2_X1 _29020_ (.A1(_05511_),
    .A2(_05562_),
    .ZN(_05563_));
 BUF_X4 _29021_ (.A(_05553_),
    .Z(_05564_));
 NAND3_X1 _29022_ (.A1(_05511_),
    .A2(_05537_),
    .A3(_05564_),
    .ZN(_05565_));
 INV_X1 _29023_ (.A(_22371_),
    .ZN(_05566_));
 INV_X1 _29024_ (.A(_22388_),
    .ZN(_05567_));
 OAI21_X1 _29025_ (.A(_05566_),
    .B1(_05567_),
    .B2(_05521_),
    .ZN(_05568_));
 INV_X1 _29026_ (.A(_22381_),
    .ZN(_05569_));
 INV_X1 _29027_ (.A(_22382_),
    .ZN(_05570_));
 AOI21_X1 _29028_ (.A(_22332_),
    .B1(_14185_),
    .B2(_22333_),
    .ZN(_05571_));
 OAI21_X2 _29029_ (.A(_05569_),
    .B1(_05570_),
    .B2(_05571_),
    .ZN(_05572_));
 OR2_X1 _29030_ (.A1(_05527_),
    .A2(_05518_),
    .ZN(_05573_));
 AOI21_X1 _29031_ (.A(_05573_),
    .B1(_05566_),
    .B2(_05521_),
    .ZN(_05574_));
 AOI221_X2 _29032_ (.A(_22364_),
    .B1(_05528_),
    .B2(_05568_),
    .C1(_05572_),
    .C2(_05574_),
    .ZN(_05575_));
 INV_X1 _29033_ (.A(_05526_),
    .ZN(_05576_));
 OAI21_X1 _29034_ (.A(_05545_),
    .B1(_05575_),
    .B2(_05576_),
    .ZN(_05577_));
 OAI21_X1 _29035_ (.A(_05512_),
    .B1(_05524_),
    .B2(_22375_),
    .ZN(_05578_));
 INV_X1 _29036_ (.A(_05578_),
    .ZN(_05579_));
 AND2_X1 _29037_ (.A1(_05577_),
    .A2(_05579_),
    .ZN(_05580_));
 OR2_X1 _29038_ (.A1(_05511_),
    .A2(_05562_),
    .ZN(_05581_));
 NAND2_X1 _29039_ (.A1(_05537_),
    .A2(_05564_),
    .ZN(_05582_));
 AOI21_X2 _29040_ (.A(_05582_),
    .B1(_05579_),
    .B2(_05577_),
    .ZN(_05583_));
 OAI221_X1 _29041_ (.A(_05563_),
    .B1(_05565_),
    .B2(_05580_),
    .C1(_05581_),
    .C2(_05583_),
    .ZN(_05584_));
 NAND4_X2 _29042_ (.A1(_05512_),
    .A2(_05564_),
    .A3(_05540_),
    .A4(_05546_),
    .ZN(_05585_));
 NOR2_X1 _29043_ (.A1(_05512_),
    .A2(_05510_),
    .ZN(_05586_));
 AND3_X1 _29044_ (.A1(_05542_),
    .A2(_05544_),
    .A3(_05545_),
    .ZN(_05587_));
 INV_X1 _29045_ (.A(_05540_),
    .ZN(_05588_));
 OAI21_X2 _29046_ (.A(_05586_),
    .B1(_05587_),
    .B2(_05588_),
    .ZN(_05589_));
 OR4_X2 _29047_ (.A1(_05512_),
    .A2(_05553_),
    .A3(_05522_),
    .A4(_05531_),
    .ZN(_05590_));
 AND2_X1 _29048_ (.A1(_05512_),
    .A2(_05510_),
    .ZN(_05591_));
 OAI21_X2 _29049_ (.A(_05591_),
    .B1(_05531_),
    .B2(_05522_),
    .ZN(_05592_));
 NAND4_X4 _29050_ (.A1(_05585_),
    .A2(_05589_),
    .A3(_05590_),
    .A4(_05592_),
    .ZN(_05593_));
 OR2_X1 _29051_ (.A1(_05553_),
    .A2(_05561_),
    .ZN(_05594_));
 NOR2_X1 _29052_ (.A1(_22354_),
    .A2(_05510_),
    .ZN(_05595_));
 OAI21_X2 _29053_ (.A(_05595_),
    .B1(_05575_),
    .B2(_05576_),
    .ZN(_05596_));
 AND3_X2 _29054_ (.A1(_05524_),
    .A2(_05594_),
    .A3(_05596_),
    .ZN(_05597_));
 AOI21_X4 _29055_ (.A(_05524_),
    .B1(_05594_),
    .B2(_05596_),
    .ZN(_05598_));
 NOR2_X4 _29056_ (.A1(_05597_),
    .A2(_05598_),
    .ZN(_05599_));
 AOI21_X1 _29057_ (.A(_05518_),
    .B1(_05566_),
    .B2(_05521_),
    .ZN(_05600_));
 AOI21_X1 _29058_ (.A(_05568_),
    .B1(_05572_),
    .B2(_05600_),
    .ZN(_05601_));
 INV_X1 _29059_ (.A(_22368_),
    .ZN(_05602_));
 OAI221_X1 _29060_ (.A(_05602_),
    .B1(_05556_),
    .B2(_05557_),
    .C1(_05558_),
    .C2(_05559_),
    .ZN(_05603_));
 MUX2_X2 _29061_ (.A(_05601_),
    .B(_05603_),
    .S(_05510_),
    .Z(_05604_));
 XNOR2_X2 _29062_ (.A(_05527_),
    .B(_05604_),
    .ZN(_05605_));
 NOR2_X1 _29063_ (.A1(_05553_),
    .A2(_05520_),
    .ZN(_05606_));
 OAI21_X2 _29064_ (.A(_05567_),
    .B1(_05541_),
    .B2(_05518_),
    .ZN(_05607_));
 AOI21_X4 _29065_ (.A(_05606_),
    .B1(_05607_),
    .B2(_05553_),
    .ZN(_05608_));
 XNOR2_X2 _29066_ (.A(_05559_),
    .B(_05608_),
    .ZN(_05609_));
 AND2_X1 _29067_ (.A1(_05553_),
    .A2(_05572_),
    .ZN(_05610_));
 INV_X1 _29068_ (.A(_05516_),
    .ZN(_05611_));
 NOR2_X1 _29069_ (.A1(_05611_),
    .A2(_05556_),
    .ZN(_05612_));
 NOR3_X1 _29070_ (.A1(_22336_),
    .A2(_05553_),
    .A3(_05612_),
    .ZN(_05613_));
 OR3_X1 _29071_ (.A1(_05519_),
    .A2(_05610_),
    .A3(_05613_),
    .ZN(_05614_));
 OAI21_X1 _29072_ (.A(_05519_),
    .B1(_05610_),
    .B2(_05613_),
    .ZN(_05615_));
 XOR2_X1 _29073_ (.A(_14183_),
    .B(_05516_),
    .Z(_05616_));
 XOR2_X1 _29074_ (.A(_14187_),
    .B(_22382_),
    .Z(_05617_));
 MUX2_X2 _29075_ (.A(_05616_),
    .B(_05617_),
    .S(_05553_),
    .Z(_05618_));
 INV_X2 _29076_ (.A(_05618_),
    .ZN(_05619_));
 AND2_X1 _29077_ (.A1(_14184_),
    .A2(_05509_),
    .ZN(_05620_));
 AOI21_X4 _29078_ (.A(_05620_),
    .B1(_05564_),
    .B2(_14188_),
    .ZN(_05621_));
 AOI22_X2 _29079_ (.A1(_05614_),
    .A2(_05615_),
    .B1(_05619_),
    .B2(_05621_),
    .ZN(_05622_));
 OAI21_X2 _29080_ (.A(_05605_),
    .B1(_05609_),
    .B2(_05622_),
    .ZN(_05623_));
 AND4_X2 _29081_ (.A1(_05585_),
    .A2(_05589_),
    .A3(_05590_),
    .A4(_05592_),
    .ZN(_05624_));
 NAND3_X2 _29082_ (.A1(_05564_),
    .A2(_05542_),
    .A3(_05544_),
    .ZN(_05625_));
 NAND2_X1 _29083_ (.A1(_22361_),
    .A2(_05510_),
    .ZN(_05626_));
 NAND2_X1 _29084_ (.A1(_05527_),
    .A2(_05510_),
    .ZN(_05627_));
 AOI21_X2 _29085_ (.A(_22368_),
    .B1(_05520_),
    .B2(_05521_),
    .ZN(_05628_));
 OAI211_X4 _29086_ (.A(_05625_),
    .B(_05626_),
    .C1(_05627_),
    .C2(_05628_),
    .ZN(_05629_));
 XNOR2_X2 _29087_ (.A(_05526_),
    .B(_05629_),
    .ZN(_05630_));
 NOR2_X1 _29088_ (.A1(_05624_),
    .A2(_05630_),
    .ZN(_05631_));
 AOI221_X1 _29089_ (.A(_05584_),
    .B1(_05593_),
    .B2(_05599_),
    .C1(_05623_),
    .C2(_05631_),
    .ZN(_05632_));
 CLKBUF_X3 _29090_ (.A(_05632_),
    .Z(_05633_));
 NOR2_X1 _29091_ (.A1(_05550_),
    .A2(_05633_),
    .ZN(_05634_));
 BUF_X4 _29092_ (.A(_05510_),
    .Z(_05635_));
 OR2_X1 _29093_ (.A1(_22340_),
    .A2(_05580_),
    .ZN(_05636_));
 AOI21_X2 _29094_ (.A(_22347_),
    .B1(_05636_),
    .B2(_05511_),
    .ZN(_05637_));
 OR2_X2 _29095_ (.A1(_05635_),
    .A2(_05637_),
    .ZN(_05638_));
 NOR2_X1 _29096_ (.A1(_05634_),
    .A2(_05638_),
    .ZN(_05639_));
 AND2_X1 _29097_ (.A1(_05535_),
    .A2(_05549_),
    .ZN(_05640_));
 CLKBUF_X3 _29098_ (.A(_05640_),
    .Z(_05641_));
 NOR2_X1 _29099_ (.A1(_05641_),
    .A2(_05633_),
    .ZN(_05642_));
 NOR3_X1 _29100_ (.A1(_05512_),
    .A2(_05524_),
    .A3(_05561_),
    .ZN(_05643_));
 NOR3_X2 _29101_ (.A1(_22343_),
    .A2(_05643_),
    .A3(_05551_),
    .ZN(_05644_));
 NOR2_X1 _29102_ (.A1(_05511_),
    .A2(_05644_),
    .ZN(_05645_));
 NOR2_X2 _29103_ (.A1(_22350_),
    .A2(_05645_),
    .ZN(_05646_));
 NOR2_X2 _29104_ (.A1(_05564_),
    .A2(_05646_),
    .ZN(_05647_));
 NOR2_X1 _29105_ (.A1(_05642_),
    .A2(_05647_),
    .ZN(_05648_));
 INV_X1 _29106_ (.A(_05490_),
    .ZN(_05649_));
 AOI21_X2 _29107_ (.A(_05649_),
    .B1(_05427_),
    .B2(_05423_),
    .ZN(_05650_));
 OAI221_X2 _29108_ (.A(_05650_),
    .B1(_05449_),
    .B2(_05443_),
    .C1(_05384_),
    .C2(_05389_),
    .ZN(_05651_));
 BUF_X4 _29109_ (.A(_05651_),
    .Z(_05652_));
 MUX2_X2 _29110_ (.A(_05639_),
    .B(_05648_),
    .S(_05652_),
    .Z(_05653_));
 OAI211_X2 _29111_ (.A(_05423_),
    .B(_05427_),
    .C1(_05498_),
    .C2(_05499_),
    .ZN(_05654_));
 INV_X1 _29112_ (.A(_05476_),
    .ZN(_05655_));
 OAI222_X2 _29113_ (.A1(_05486_),
    .A2(_05483_),
    .B1(_05416_),
    .B2(_05655_),
    .C1(_05467_),
    .C2(_05411_),
    .ZN(_05656_));
 AOI221_X1 _29114_ (.A(_05564_),
    .B1(_05654_),
    .B2(_05656_),
    .C1(_05471_),
    .C2(_05470_),
    .ZN(_05657_));
 AND2_X1 _29115_ (.A1(_05487_),
    .A2(_05635_),
    .ZN(_05658_));
 AOI221_X4 _29116_ (.A(_05657_),
    .B1(_05658_),
    .B2(_05390_),
    .C1(_05400_),
    .C2(_05635_),
    .ZN(_05659_));
 AOI22_X2 _29117_ (.A1(_05470_),
    .A2(_05471_),
    .B1(_05654_),
    .B2(_05656_),
    .ZN(_05660_));
 AND3_X1 _29118_ (.A1(_05470_),
    .A2(_05471_),
    .A3(_05487_),
    .ZN(_05661_));
 OR4_X4 _29119_ (.A1(_05400_),
    .A2(_05635_),
    .A3(_05660_),
    .A4(_05661_),
    .ZN(_05662_));
 NAND2_X2 _29120_ (.A1(_05641_),
    .A2(_05652_),
    .ZN(_05663_));
 MUX2_X2 _29121_ (.A(_22392_),
    .B(_22394_),
    .S(_05564_),
    .Z(_05664_));
 NOR2_X1 _29122_ (.A1(_05618_),
    .A2(_05664_),
    .ZN(_05665_));
 INV_X1 _29123_ (.A(_05665_),
    .ZN(_05666_));
 AOI21_X1 _29124_ (.A(_05630_),
    .B1(_05609_),
    .B2(_05605_),
    .ZN(_05667_));
 OAI21_X2 _29125_ (.A(_05593_),
    .B1(_05599_),
    .B2(_05667_),
    .ZN(_05668_));
 NOR2_X1 _29126_ (.A1(_05562_),
    .A2(_05583_),
    .ZN(_05669_));
 XNOR2_X2 _29127_ (.A(_05511_),
    .B(_05669_),
    .ZN(_05670_));
 AOI221_X2 _29128_ (.A(_05502_),
    .B1(_05503_),
    .B2(_05504_),
    .C1(_05470_),
    .C2(_05471_),
    .ZN(_05671_));
 BUF_X4 _29129_ (.A(_05671_),
    .Z(_05672_));
 AOI221_X2 _29130_ (.A(_05666_),
    .B1(_05668_),
    .B2(_05670_),
    .C1(_05672_),
    .C2(_05550_),
    .ZN(_05673_));
 NAND4_X4 _29131_ (.A1(_05659_),
    .A2(_05662_),
    .A3(_05663_),
    .A4(_05673_),
    .ZN(_05674_));
 NAND2_X2 _29132_ (.A1(_05653_),
    .A2(_05674_),
    .ZN(_22396_));
 INV_X1 _29133_ (.A(_22396_),
    .ZN(_22398_));
 OAI21_X2 _29134_ (.A(_05650_),
    .B1(_05449_),
    .B2(_05443_),
    .ZN(_05675_));
 BUF_X1 _29135_ (.A(_22401_),
    .Z(_05676_));
 INV_X1 _29136_ (.A(_05676_),
    .ZN(_05677_));
 AOI21_X1 _29137_ (.A(_22347_),
    .B1(_05548_),
    .B2(_05636_),
    .ZN(_05678_));
 OR2_X1 _29138_ (.A1(_05510_),
    .A2(_05678_),
    .ZN(_05679_));
 NAND2_X1 _29139_ (.A1(_05677_),
    .A2(_05679_),
    .ZN(_05680_));
 XNOR2_X2 _29140_ (.A(_05528_),
    .B(_05604_),
    .ZN(_05681_));
 AND2_X1 _29141_ (.A1(_05614_),
    .A2(_05615_),
    .ZN(_05682_));
 BUF_X2 _29142_ (.A(_05682_),
    .Z(_05683_));
 NOR4_X1 _29143_ (.A1(_05681_),
    .A2(_05609_),
    .A3(_05683_),
    .A4(_05618_),
    .ZN(_05684_));
 XNOR2_X2 _29144_ (.A(_05576_),
    .B(_05629_),
    .ZN(_05685_));
 OAI211_X4 _29145_ (.A(_05593_),
    .B(_05685_),
    .C1(_05598_),
    .C2(_05597_),
    .ZN(_05686_));
 OR3_X2 _29146_ (.A1(_05584_),
    .A2(_05684_),
    .A3(_05686_),
    .ZN(_05687_));
 NOR2_X1 _29147_ (.A1(_05635_),
    .A2(_05678_),
    .ZN(_05688_));
 NAND3_X1 _29148_ (.A1(_05676_),
    .A2(_05687_),
    .A3(_05688_),
    .ZN(_05689_));
 AOI221_X1 _29149_ (.A(_05675_),
    .B1(_05680_),
    .B2(_05689_),
    .C1(_05471_),
    .C2(_05470_),
    .ZN(_05690_));
 INV_X1 _29150_ (.A(_22350_),
    .ZN(_05691_));
 OAI21_X2 _29151_ (.A(_05691_),
    .B1(_05511_),
    .B2(_05644_),
    .ZN(_05692_));
 OAI21_X2 _29152_ (.A(_05549_),
    .B1(_05692_),
    .B2(_05535_),
    .ZN(_05693_));
 NAND2_X1 _29153_ (.A1(_05687_),
    .A2(_05693_),
    .ZN(_05694_));
 AOI211_X2 _29154_ (.A(_05677_),
    .B(_05694_),
    .C1(_05505_),
    .C2(_05472_),
    .ZN(_05695_));
 OR2_X1 _29155_ (.A1(_05676_),
    .A2(_05693_),
    .ZN(_05696_));
 OR3_X1 _29156_ (.A1(_05384_),
    .A2(_05389_),
    .A3(_05696_),
    .ZN(_05697_));
 OAI221_X1 _29157_ (.A(_05697_),
    .B1(_05696_),
    .B2(_05505_),
    .C1(_05676_),
    .C2(_05687_),
    .ZN(_05698_));
 OR3_X2 _29158_ (.A1(_05690_),
    .A2(_05695_),
    .A3(_05698_),
    .ZN(_05699_));
 INV_X2 _29159_ (.A(_05699_),
    .ZN(_22422_));
 MUX2_X2 _29160_ (.A(_05688_),
    .B(_05693_),
    .S(_05652_),
    .Z(_05700_));
 CLKBUF_X3 _29161_ (.A(_05700_),
    .Z(_05701_));
 CLKBUF_X3 _29162_ (.A(_14190_),
    .Z(_05702_));
 INV_X2 _29163_ (.A(_05702_),
    .ZN(_05703_));
 AOI221_X1 _29164_ (.A(_05703_),
    .B1(_05672_),
    .B2(_05638_),
    .C1(_05692_),
    .C2(_05635_),
    .ZN(_05704_));
 NOR4_X4 _29165_ (.A1(_05584_),
    .A2(_05681_),
    .A3(_05609_),
    .A4(_05686_),
    .ZN(_05705_));
 OR2_X1 _29166_ (.A1(_05683_),
    .A2(_05618_),
    .ZN(_05706_));
 NAND2_X1 _29167_ (.A1(_05593_),
    .A2(_05706_),
    .ZN(_05707_));
 AOI21_X4 _29168_ (.A(_05599_),
    .B1(_05623_),
    .B2(_05685_),
    .ZN(_05708_));
 OAI21_X2 _29169_ (.A(_05705_),
    .B1(_05707_),
    .B2(_05708_),
    .ZN(_05709_));
 XNOR2_X1 _29170_ (.A(_05677_),
    .B(_05687_),
    .ZN(_05710_));
 AND2_X1 _29171_ (.A1(_05709_),
    .A2(_05710_),
    .ZN(_05711_));
 NAND3_X1 _29172_ (.A1(_05701_),
    .A2(_05704_),
    .A3(_05711_),
    .ZN(_05712_));
 CLKBUF_X2 _29173_ (.A(_22397_),
    .Z(_05713_));
 CLKBUF_X3 _29174_ (.A(_05713_),
    .Z(_05714_));
 NAND3_X1 _29175_ (.A1(_05714_),
    .A2(_05621_),
    .A3(_05664_),
    .ZN(_05715_));
 BUF_X4 _29176_ (.A(_05701_),
    .Z(_05716_));
 OAI21_X1 _29177_ (.A(_05712_),
    .B1(_05715_),
    .B2(_05716_),
    .ZN(_05717_));
 NAND2_X2 _29178_ (.A1(_05659_),
    .A2(_05662_),
    .ZN(_05718_));
 AND2_X1 _29179_ (.A1(_22392_),
    .A2(_05635_),
    .ZN(_05719_));
 AOI21_X4 _29180_ (.A(_05719_),
    .B1(_05564_),
    .B2(_22394_),
    .ZN(_05720_));
 NOR4_X1 _29181_ (.A1(_05714_),
    .A2(_05718_),
    .A3(_05720_),
    .A4(_05701_),
    .ZN(_05721_));
 XNOR2_X2 _29182_ (.A(_05550_),
    .B(_05672_),
    .ZN(_05722_));
 OAI21_X1 _29183_ (.A(_05633_),
    .B1(_05666_),
    .B2(_05668_),
    .ZN(_05723_));
 NAND2_X1 _29184_ (.A1(_05704_),
    .A2(_05723_),
    .ZN(_05724_));
 NOR2_X1 _29185_ (.A1(_05703_),
    .A2(_05664_),
    .ZN(_05725_));
 AND4_X2 _29186_ (.A1(_05659_),
    .A2(_05662_),
    .A3(_05663_),
    .A4(_05673_),
    .ZN(_05726_));
 OR2_X1 _29187_ (.A1(_05634_),
    .A2(_05638_),
    .ZN(_05727_));
 NAND2_X2 _29188_ (.A1(_05635_),
    .A2(_05692_),
    .ZN(_05728_));
 OAI21_X1 _29189_ (.A(_05728_),
    .B1(_05633_),
    .B2(_05641_),
    .ZN(_05729_));
 MUX2_X1 _29190_ (.A(_05727_),
    .B(_05729_),
    .S(_05652_),
    .Z(_05730_));
 OAI33_X1 _29191_ (.A1(_05718_),
    .A2(_05722_),
    .A3(_05724_),
    .B1(_05725_),
    .B2(_05726_),
    .B3(_05730_),
    .ZN(_05731_));
 INV_X1 _29192_ (.A(_05713_),
    .ZN(_05732_));
 BUF_X4 _29193_ (.A(_05732_),
    .Z(_05733_));
 AOI21_X2 _29194_ (.A(_05701_),
    .B1(_05720_),
    .B2(_05733_),
    .ZN(_05734_));
 OAI21_X4 _29195_ (.A(_05670_),
    .B1(_05624_),
    .B2(_05708_),
    .ZN(_05735_));
 XNOR2_X2 _29196_ (.A(_05641_),
    .B(_05672_),
    .ZN(_05736_));
 NAND2_X4 _29197_ (.A1(_05735_),
    .A2(_05736_),
    .ZN(_05737_));
 CLKBUF_X3 _29198_ (.A(_05736_),
    .Z(_05738_));
 NAND3_X1 _29199_ (.A1(_05735_),
    .A2(_05738_),
    .A3(_05704_),
    .ZN(_05739_));
 AOI22_X2 _29200_ (.A1(_05701_),
    .A2(_05737_),
    .B1(_05739_),
    .B2(_05733_),
    .ZN(_05740_));
 AND2_X2 _29201_ (.A1(_05659_),
    .A2(_05662_),
    .ZN(_05741_));
 OAI222_X2 _29202_ (.A1(_05717_),
    .A2(_05721_),
    .B1(_05731_),
    .B2(_05734_),
    .C1(_05740_),
    .C2(_05741_),
    .ZN(_05742_));
 INV_X1 _29203_ (.A(_05742_),
    .ZN(_22403_));
 INV_X1 _29204_ (.A(_05693_),
    .ZN(_05743_));
 MUX2_X1 _29205_ (.A(_05679_),
    .B(_05743_),
    .S(_05652_),
    .Z(_05744_));
 CLKBUF_X3 _29206_ (.A(_05744_),
    .Z(_05745_));
 BUF_X4 _29207_ (.A(_05745_),
    .Z(_05746_));
 OAI21_X1 _29208_ (.A(_05746_),
    .B1(_05741_),
    .B2(_05714_),
    .ZN(_05747_));
 NAND2_X1 _29209_ (.A1(_05701_),
    .A2(_05711_),
    .ZN(_05748_));
 CLKBUF_X3 _29210_ (.A(_05702_),
    .Z(_05749_));
 AOI21_X4 _29211_ (.A(_05647_),
    .B1(_05638_),
    .B2(_05672_),
    .ZN(_05750_));
 NAND2_X1 _29212_ (.A1(_05749_),
    .A2(_05750_),
    .ZN(_05751_));
 AOI22_X1 _29213_ (.A1(_05659_),
    .A2(_05662_),
    .B1(_05738_),
    .B2(_05735_),
    .ZN(_05752_));
 OR2_X1 _29214_ (.A1(_05751_),
    .A2(_05752_),
    .ZN(_05753_));
 OAI21_X1 _29215_ (.A(_05747_),
    .B1(_05748_),
    .B2(_05753_),
    .ZN(_05754_));
 NOR2_X2 _29216_ (.A1(_05733_),
    .A2(_05701_),
    .ZN(_05755_));
 NAND2_X1 _29217_ (.A1(_05720_),
    .A2(_05755_),
    .ZN(_05756_));
 NAND2_X1 _29218_ (.A1(_05754_),
    .A2(_05756_),
    .ZN(_05757_));
 BUF_X4 _29219_ (.A(_05699_),
    .Z(_05758_));
 NOR2_X2 _29220_ (.A1(_05635_),
    .A2(_05637_),
    .ZN(_05759_));
 OAI21_X4 _29221_ (.A(_05728_),
    .B1(_05759_),
    .B2(_05652_),
    .ZN(_05760_));
 NOR2_X1 _29222_ (.A1(_05679_),
    .A2(_05709_),
    .ZN(_05761_));
 NOR2_X1 _29223_ (.A1(_05743_),
    .A2(_05709_),
    .ZN(_05762_));
 MUX2_X1 _29224_ (.A(_05761_),
    .B(_05762_),
    .S(_05652_),
    .Z(_05763_));
 OR2_X1 _29225_ (.A1(_05760_),
    .A2(_05763_),
    .ZN(_05764_));
 BUF_X4 _29226_ (.A(_05764_),
    .Z(_05765_));
 NOR2_X1 _29227_ (.A1(_05758_),
    .A2(_05765_),
    .ZN(_05766_));
 AOI21_X1 _29228_ (.A(_05746_),
    .B1(_05766_),
    .B2(_22399_),
    .ZN(_05767_));
 NOR2_X1 _29229_ (.A1(_05757_),
    .A2(_05767_),
    .ZN(_05768_));
 AND2_X2 _29230_ (.A1(_05700_),
    .A2(_05711_),
    .ZN(_05769_));
 AOI21_X1 _29231_ (.A(_05734_),
    .B1(_05769_),
    .B2(_05731_),
    .ZN(_05770_));
 MUX2_X2 _29232_ (.A(_14188_),
    .B(_14184_),
    .S(_05635_),
    .Z(_05771_));
 AOI21_X1 _29233_ (.A(_05770_),
    .B1(_05755_),
    .B2(_05771_),
    .ZN(_05772_));
 MUX2_X1 _29234_ (.A(_05768_),
    .B(_05757_),
    .S(_05772_),
    .Z(_05773_));
 BUF_X4 _29235_ (.A(_05703_),
    .Z(_05774_));
 AOI21_X2 _29236_ (.A(_05605_),
    .B1(_05735_),
    .B2(_05738_),
    .ZN(_05775_));
 XNOR2_X2 _29237_ (.A(_05521_),
    .B(_05608_),
    .ZN(_05776_));
 NOR3_X1 _29238_ (.A1(_05776_),
    .A2(_05633_),
    .A3(_05722_),
    .ZN(_05777_));
 OAI21_X2 _29239_ (.A(_05774_),
    .B1(_05775_),
    .B2(_05777_),
    .ZN(_05778_));
 OAI21_X1 _29240_ (.A(_05685_),
    .B1(_05593_),
    .B2(_05584_),
    .ZN(_05779_));
 NOR2_X1 _29241_ (.A1(_05641_),
    .A2(_05779_),
    .ZN(_05780_));
 OR2_X1 _29242_ (.A1(_05550_),
    .A2(_05779_),
    .ZN(_05781_));
 AOI21_X1 _29243_ (.A(_05781_),
    .B1(_05471_),
    .B2(_05470_),
    .ZN(_05782_));
 MUX2_X1 _29244_ (.A(_05780_),
    .B(_05782_),
    .S(_05505_),
    .Z(_05783_));
 NOR4_X2 _29245_ (.A1(_05390_),
    .A2(_05675_),
    .A3(_05641_),
    .A4(_05599_),
    .ZN(_05784_));
 OR2_X1 _29246_ (.A1(_05550_),
    .A2(_05599_),
    .ZN(_05785_));
 NOR2_X1 _29247_ (.A1(_05505_),
    .A2(_05785_),
    .ZN(_05786_));
 NAND3_X1 _29248_ (.A1(_05470_),
    .A2(_05471_),
    .A3(_05780_),
    .ZN(_05787_));
 OAI221_X2 _29249_ (.A(_05787_),
    .B1(_05599_),
    .B2(_05584_),
    .C1(_05472_),
    .C2(_05785_),
    .ZN(_05788_));
 NOR4_X2 _29250_ (.A1(_05783_),
    .A2(_05784_),
    .A3(_05786_),
    .A4(_05788_),
    .ZN(_05789_));
 AOI21_X2 _29251_ (.A(_05765_),
    .B1(_05789_),
    .B2(_05749_),
    .ZN(_05790_));
 AOI22_X2 _29252_ (.A1(_05778_),
    .A2(_05790_),
    .B1(_05753_),
    .B2(_05765_),
    .ZN(_05791_));
 NOR2_X1 _29253_ (.A1(_22422_),
    .A2(_05791_),
    .ZN(_05792_));
 NOR2_X1 _29254_ (.A1(_05702_),
    .A2(_05771_),
    .ZN(_05793_));
 AOI21_X1 _29255_ (.A(_05793_),
    .B1(_05683_),
    .B2(_05702_),
    .ZN(_05794_));
 NOR2_X1 _29256_ (.A1(_05760_),
    .A2(_05794_),
    .ZN(_05795_));
 NAND3_X1 _29257_ (.A1(_05674_),
    .A2(_05737_),
    .A3(_05795_),
    .ZN(_05796_));
 MUX2_X1 _29258_ (.A(_05618_),
    .B(_05664_),
    .S(_05703_),
    .Z(_05797_));
 OAI221_X2 _29259_ (.A(_05797_),
    .B1(_05759_),
    .B2(_05652_),
    .C1(_05564_),
    .C2(_05646_),
    .ZN(_05798_));
 NOR2_X4 _29260_ (.A1(_05633_),
    .A2(_05722_),
    .ZN(_05799_));
 NOR2_X1 _29261_ (.A1(_05726_),
    .A2(_05799_),
    .ZN(_05800_));
 OAI21_X2 _29262_ (.A(_05796_),
    .B1(_05798_),
    .B2(_05800_),
    .ZN(_05801_));
 AOI21_X2 _29263_ (.A(_05670_),
    .B1(_05593_),
    .B2(_05738_),
    .ZN(_05802_));
 AOI221_X2 _29264_ (.A(_05758_),
    .B1(_05765_),
    .B2(_05801_),
    .C1(_05802_),
    .C2(_05774_),
    .ZN(_05803_));
 NOR3_X2 _29265_ (.A1(_05746_),
    .A2(_05792_),
    .A3(_05803_),
    .ZN(_05804_));
 AOI21_X4 _29266_ (.A(_05804_),
    .B1(_05760_),
    .B2(_05733_),
    .ZN(_05805_));
 AOI21_X1 _29267_ (.A(_22399_),
    .B1(_05750_),
    .B2(_05709_),
    .ZN(_05806_));
 OR2_X1 _29268_ (.A1(_05745_),
    .A2(_05806_),
    .ZN(_05807_));
 MUX2_X1 _29269_ (.A(_05681_),
    .B(_05630_),
    .S(_05653_),
    .Z(_05808_));
 INV_X1 _29270_ (.A(_05808_),
    .ZN(_05809_));
 NOR3_X1 _29271_ (.A1(_05774_),
    .A2(_05699_),
    .A3(_05765_),
    .ZN(_05810_));
 NAND2_X1 _29272_ (.A1(_05670_),
    .A2(_05668_),
    .ZN(_05811_));
 AND3_X1 _29273_ (.A1(_05683_),
    .A2(_05811_),
    .A3(_05738_),
    .ZN(_05812_));
 NOR3_X1 _29274_ (.A1(_05702_),
    .A2(_05641_),
    .A3(_05633_),
    .ZN(_05813_));
 OR3_X1 _29275_ (.A1(_05702_),
    .A2(_05550_),
    .A3(_05633_),
    .ZN(_05814_));
 AOI21_X1 _29276_ (.A(_05814_),
    .B1(_05471_),
    .B2(_05470_),
    .ZN(_05815_));
 MUX2_X1 _29277_ (.A(_05813_),
    .B(_05815_),
    .S(_05505_),
    .Z(_05816_));
 AOI221_X2 _29278_ (.A(_05816_),
    .B1(_05813_),
    .B2(_05390_),
    .C1(_05703_),
    .C2(_05776_),
    .ZN(_05817_));
 OAI21_X1 _29279_ (.A(_05750_),
    .B1(_05812_),
    .B2(_05817_),
    .ZN(_05818_));
 AOI221_X2 _29280_ (.A(_05807_),
    .B1(_05809_),
    .B2(_05810_),
    .C1(_05818_),
    .C2(_05766_),
    .ZN(_05819_));
 NAND2_X1 _29281_ (.A1(_05702_),
    .A2(_05771_),
    .ZN(_05820_));
 AND2_X1 _29282_ (.A1(_05750_),
    .A2(_05820_),
    .ZN(_05821_));
 OAI221_X2 _29283_ (.A(_05821_),
    .B1(_05799_),
    .B2(_05726_),
    .C1(_05749_),
    .C2(_05741_),
    .ZN(_05822_));
 AOI21_X1 _29284_ (.A(_05798_),
    .B1(_05738_),
    .B2(_05735_),
    .ZN(_05823_));
 NOR2_X1 _29285_ (.A1(_22422_),
    .A2(_05823_),
    .ZN(_05824_));
 AOI22_X4 _29286_ (.A1(_05758_),
    .A2(_05765_),
    .B1(_05822_),
    .B2(_05824_),
    .ZN(_05825_));
 MUX2_X1 _29287_ (.A(_05599_),
    .B(_05630_),
    .S(_05733_),
    .Z(_05826_));
 AOI22_X4 _29288_ (.A1(_05819_),
    .A2(_05825_),
    .B1(_05826_),
    .B2(_05746_),
    .ZN(_05827_));
 OR2_X1 _29289_ (.A1(_05708_),
    .A2(_05707_),
    .ZN(_05828_));
 AOI21_X2 _29290_ (.A(_05710_),
    .B1(_05828_),
    .B2(_05705_),
    .ZN(_05829_));
 AND2_X1 _29291_ (.A1(_05716_),
    .A2(_05829_),
    .ZN(_05830_));
 NAND2_X1 _29292_ (.A1(_05701_),
    .A2(_22422_),
    .ZN(_05831_));
 AOI221_X2 _29293_ (.A(_05831_),
    .B1(_05790_),
    .B2(_05778_),
    .C1(_05765_),
    .C2(_05753_),
    .ZN(_05832_));
 MUX2_X1 _29294_ (.A(_05624_),
    .B(_05599_),
    .S(_05733_),
    .Z(_05833_));
 AOI222_X2 _29295_ (.A1(_05801_),
    .A2(_05830_),
    .B1(_05832_),
    .B2(_05819_),
    .C1(_05833_),
    .C2(_05745_),
    .ZN(_05834_));
 MUX2_X1 _29296_ (.A(_05584_),
    .B(_05624_),
    .S(_05733_),
    .Z(_05835_));
 NOR2_X1 _29297_ (.A1(_05716_),
    .A2(_05835_),
    .ZN(_05836_));
 INV_X1 _29298_ (.A(_05765_),
    .ZN(_22426_));
 NAND2_X1 _29299_ (.A1(_22422_),
    .A2(_22426_),
    .ZN(_05837_));
 OAI211_X2 _29300_ (.A(_05624_),
    .B(_05750_),
    .C1(_05722_),
    .C2(_05670_),
    .ZN(_05838_));
 NAND2_X1 _29301_ (.A1(_05550_),
    .A2(_05672_),
    .ZN(_05839_));
 NAND2_X1 _29302_ (.A1(_05641_),
    .A2(_05728_),
    .ZN(_05840_));
 OAI221_X2 _29303_ (.A(_05599_),
    .B1(_05638_),
    .B2(_05839_),
    .C1(_05840_),
    .C2(_05672_),
    .ZN(_05841_));
 AND3_X1 _29304_ (.A1(_05749_),
    .A2(_05838_),
    .A3(_05841_),
    .ZN(_05842_));
 NOR2_X1 _29305_ (.A1(_05749_),
    .A2(_05808_),
    .ZN(_05843_));
 OAI211_X2 _29306_ (.A(_05774_),
    .B(_05771_),
    .C1(_05730_),
    .C2(_05619_),
    .ZN(_05844_));
 NOR2_X1 _29307_ (.A1(_05702_),
    .A2(_05618_),
    .ZN(_05845_));
 NAND2_X1 _29308_ (.A1(_05653_),
    .A2(_05845_),
    .ZN(_05846_));
 OAI21_X1 _29309_ (.A(_05844_),
    .B1(_05846_),
    .B2(_05726_),
    .ZN(_05847_));
 NAND2_X1 _29310_ (.A1(_05758_),
    .A2(_22426_),
    .ZN(_05848_));
 NAND3_X1 _29311_ (.A1(_05683_),
    .A2(_05811_),
    .A3(_05738_),
    .ZN(_05849_));
 AOI21_X1 _29312_ (.A(_05774_),
    .B1(_05609_),
    .B2(_05653_),
    .ZN(_05850_));
 AND2_X1 _29313_ (.A1(_05849_),
    .A2(_05850_),
    .ZN(_05851_));
 OAI33_X1 _29314_ (.A1(_05837_),
    .A2(_05842_),
    .A3(_05843_),
    .B1(_05847_),
    .B2(_05848_),
    .B3(_05851_),
    .ZN(_05852_));
 NOR2_X1 _29315_ (.A1(_05683_),
    .A2(_05618_),
    .ZN(_05853_));
 AND4_X1 _29316_ (.A1(_05659_),
    .A2(_05662_),
    .A3(_05704_),
    .A4(_05723_),
    .ZN(_05854_));
 NAND4_X1 _29317_ (.A1(_05677_),
    .A2(_05738_),
    .A3(_05853_),
    .A4(_05854_),
    .ZN(_05855_));
 NAND2_X1 _29318_ (.A1(_05749_),
    .A2(_05720_),
    .ZN(_05856_));
 NAND3_X1 _29319_ (.A1(_05677_),
    .A2(_05853_),
    .A3(_05856_),
    .ZN(_05857_));
 AOI21_X1 _29320_ (.A(_05856_),
    .B1(_05854_),
    .B2(_05738_),
    .ZN(_05858_));
 NAND4_X1 _29321_ (.A1(_05676_),
    .A2(_05653_),
    .A3(_05674_),
    .A4(_05706_),
    .ZN(_05859_));
 OAI221_X1 _29322_ (.A(_05855_),
    .B1(_05857_),
    .B2(_22396_),
    .C1(_05858_),
    .C2(_05859_),
    .ZN(_05860_));
 AOI211_X4 _29323_ (.A(_05745_),
    .B(_05852_),
    .C1(_05860_),
    .C2(_05705_),
    .ZN(_05861_));
 NOR4_X2 _29324_ (.A1(_05827_),
    .A2(_05834_),
    .A3(_05836_),
    .A4(_05861_),
    .ZN(_05862_));
 NOR2_X1 _29325_ (.A1(_05713_),
    .A2(_05609_),
    .ZN(_05863_));
 AOI21_X1 _29326_ (.A(_05863_),
    .B1(_05605_),
    .B2(_05714_),
    .ZN(_05864_));
 NOR2_X1 _29327_ (.A1(_05716_),
    .A2(_05864_),
    .ZN(_05865_));
 NOR2_X1 _29328_ (.A1(_05763_),
    .A2(_05865_),
    .ZN(_05866_));
 INV_X1 _29329_ (.A(_05866_),
    .ZN(_05867_));
 NOR2_X1 _29330_ (.A1(_05701_),
    .A2(_05863_),
    .ZN(_05868_));
 AOI21_X1 _29331_ (.A(_05758_),
    .B1(_05849_),
    .B2(_05850_),
    .ZN(_05869_));
 AOI211_X2 _29332_ (.A(_05702_),
    .B(_05621_),
    .C1(_05653_),
    .C2(_05618_),
    .ZN(_05870_));
 AND2_X1 _29333_ (.A1(_05653_),
    .A2(_05845_),
    .ZN(_05871_));
 AOI21_X1 _29334_ (.A(_05870_),
    .B1(_05871_),
    .B2(_05674_),
    .ZN(_05872_));
 AOI221_X2 _29335_ (.A(_05868_),
    .B1(_05869_),
    .B2(_05872_),
    .C1(_05731_),
    .C2(_05758_),
    .ZN(_05873_));
 NAND2_X1 _29336_ (.A1(_05750_),
    .A2(_05820_),
    .ZN(_05874_));
 AOI221_X2 _29337_ (.A(_05874_),
    .B1(_05737_),
    .B2(_05674_),
    .C1(_05774_),
    .C2(_05718_),
    .ZN(_05875_));
 MUX2_X1 _29338_ (.A(_05683_),
    .B(_05618_),
    .S(_05732_),
    .Z(_05876_));
 AND2_X1 _29339_ (.A1(_22399_),
    .A2(_05829_),
    .ZN(_05877_));
 MUX2_X1 _29340_ (.A(_05876_),
    .B(_05877_),
    .S(_05700_),
    .Z(_05878_));
 OR2_X1 _29341_ (.A1(_05823_),
    .A2(_05878_),
    .ZN(_05879_));
 OAI22_X4 _29342_ (.A1(_05875_),
    .A2(_05879_),
    .B1(_05769_),
    .B2(_05878_),
    .ZN(_05880_));
 NAND2_X1 _29343_ (.A1(_05700_),
    .A2(_05829_),
    .ZN(_05881_));
 NOR3_X1 _29344_ (.A1(_05751_),
    .A2(_05752_),
    .A3(_05881_),
    .ZN(_05882_));
 NOR2_X1 _29345_ (.A1(_05733_),
    .A2(_05776_),
    .ZN(_05883_));
 AOI21_X1 _29346_ (.A(_05883_),
    .B1(_05683_),
    .B2(_05733_),
    .ZN(_05884_));
 NOR2_X1 _29347_ (.A1(_05701_),
    .A2(_05884_),
    .ZN(_05885_));
 AND4_X1 _29348_ (.A1(_05674_),
    .A2(_05737_),
    .A3(_05795_),
    .A4(_05769_),
    .ZN(_05886_));
 NAND4_X1 _29349_ (.A1(_05700_),
    .A2(_05750_),
    .A3(_05711_),
    .A4(_05797_),
    .ZN(_05887_));
 AOI21_X1 _29350_ (.A(_05887_),
    .B1(_05737_),
    .B2(_05674_),
    .ZN(_05888_));
 NOR4_X2 _29351_ (.A1(_05882_),
    .A2(_05885_),
    .A3(_05886_),
    .A4(_05888_),
    .ZN(_05889_));
 OR4_X1 _29352_ (.A1(_05867_),
    .A2(_05873_),
    .A3(_05880_),
    .A4(_05889_),
    .ZN(_05890_));
 AOI21_X1 _29353_ (.A(_05856_),
    .B1(_05737_),
    .B2(_05674_),
    .ZN(_05891_));
 NOR2_X1 _29354_ (.A1(_05550_),
    .A2(_05672_),
    .ZN(_05892_));
 AOI21_X1 _29355_ (.A(_05666_),
    .B1(_05668_),
    .B2(_05670_),
    .ZN(_05893_));
 OAI21_X1 _29356_ (.A(_05893_),
    .B1(_05652_),
    .B2(_05641_),
    .ZN(_05894_));
 OAI21_X1 _29357_ (.A(_05702_),
    .B1(_05892_),
    .B2(_05894_),
    .ZN(_05895_));
 AOI221_X2 _29358_ (.A(_05799_),
    .B1(_05895_),
    .B2(_05741_),
    .C1(_05621_),
    .C2(_05749_),
    .ZN(_05896_));
 NOR3_X1 _29359_ (.A1(_05881_),
    .A2(_05891_),
    .A3(_05896_),
    .ZN(_05897_));
 MUX2_X1 _29360_ (.A(_05681_),
    .B(_05630_),
    .S(_05714_),
    .Z(_05898_));
 NOR2_X1 _29361_ (.A1(_05749_),
    .A2(_05683_),
    .ZN(_05899_));
 MUX2_X1 _29362_ (.A(_05845_),
    .B(_05899_),
    .S(_05737_),
    .Z(_05900_));
 NAND2_X1 _29363_ (.A1(_05749_),
    .A2(_05605_),
    .ZN(_05901_));
 OAI33_X1 _29364_ (.A1(_05774_),
    .A2(_05609_),
    .A3(_05775_),
    .B1(_05901_),
    .B2(_05726_),
    .B3(_05799_),
    .ZN(_05902_));
 NOR2_X1 _29365_ (.A1(_05900_),
    .A2(_05902_),
    .ZN(_05903_));
 AOI221_X2 _29366_ (.A(_05897_),
    .B1(_05898_),
    .B2(_05745_),
    .C1(_05769_),
    .C2(_05903_),
    .ZN(_05904_));
 OAI21_X2 _29367_ (.A(_05745_),
    .B1(_05621_),
    .B2(_05713_),
    .ZN(_05905_));
 AOI22_X2 _29368_ (.A1(_05619_),
    .A2(_05755_),
    .B1(_05748_),
    .B2(_05905_),
    .ZN(_05906_));
 OAI211_X2 _29369_ (.A(_05725_),
    .B(_05905_),
    .C1(_05726_),
    .C2(_05799_),
    .ZN(_05907_));
 AOI21_X1 _29370_ (.A(_05774_),
    .B1(_05663_),
    .B2(_05673_),
    .ZN(_05908_));
 OAI221_X2 _29371_ (.A(_05737_),
    .B1(_05908_),
    .B2(_05718_),
    .C1(_05771_),
    .C2(_05774_),
    .ZN(_05909_));
 INV_X1 _29372_ (.A(_05905_),
    .ZN(_05910_));
 OAI211_X2 _29373_ (.A(_05906_),
    .B(_05907_),
    .C1(_05909_),
    .C2(_05910_),
    .ZN(_05911_));
 OR2_X1 _29374_ (.A1(_05742_),
    .A2(_05911_),
    .ZN(_05912_));
 NOR3_X2 _29375_ (.A1(_05890_),
    .A2(_05904_),
    .A3(_05912_),
    .ZN(_05913_));
 NAND3_X1 _29376_ (.A1(_05774_),
    .A2(_05716_),
    .A3(_05709_),
    .ZN(_05914_));
 AOI221_X2 _29377_ (.A(_22422_),
    .B1(_05750_),
    .B2(_05812_),
    .C1(_05653_),
    .C2(_05609_),
    .ZN(_05915_));
 AND3_X1 _29378_ (.A1(_22422_),
    .A2(_05838_),
    .A3(_05841_),
    .ZN(_05916_));
 NOR3_X2 _29379_ (.A1(_05914_),
    .A2(_05915_),
    .A3(_05916_),
    .ZN(_05917_));
 NOR3_X1 _29380_ (.A1(_05584_),
    .A2(_05722_),
    .A3(_05758_),
    .ZN(_05918_));
 NOR2_X1 _29381_ (.A1(_22422_),
    .A2(_05808_),
    .ZN(_05919_));
 NAND2_X1 _29382_ (.A1(_05704_),
    .A2(_22426_),
    .ZN(_05920_));
 NOR4_X2 _29383_ (.A1(_05745_),
    .A2(_05918_),
    .A3(_05919_),
    .A4(_05920_),
    .ZN(_05921_));
 MUX2_X1 _29384_ (.A(_05722_),
    .B(_05760_),
    .S(_05713_),
    .Z(_05922_));
 OR4_X1 _29385_ (.A1(_05758_),
    .A2(_05875_),
    .A3(_05823_),
    .A4(_05922_),
    .ZN(_05923_));
 NOR2_X1 _29386_ (.A1(_05763_),
    .A2(_05922_),
    .ZN(_05924_));
 NOR3_X1 _29387_ (.A1(_22399_),
    .A2(_22422_),
    .A3(_05922_),
    .ZN(_05925_));
 NOR2_X1 _29388_ (.A1(_05924_),
    .A2(_05925_),
    .ZN(_05926_));
 AOI211_X2 _29389_ (.A(_05917_),
    .B(_05921_),
    .C1(_05923_),
    .C2(_05926_),
    .ZN(_05927_));
 MUX2_X1 _29390_ (.A(_05670_),
    .B(_05738_),
    .S(_05714_),
    .Z(_05928_));
 NOR2_X1 _29391_ (.A1(_05716_),
    .A2(_05928_),
    .ZN(_05929_));
 MUX2_X1 _29392_ (.A(_05789_),
    .B(_05802_),
    .S(_05749_),
    .Z(_05930_));
 NOR2_X1 _29393_ (.A1(_05745_),
    .A2(_05758_),
    .ZN(_05931_));
 OR3_X1 _29394_ (.A1(_05758_),
    .A2(_05760_),
    .A3(_05709_),
    .ZN(_05932_));
 OAI33_X1 _29395_ (.A1(_22422_),
    .A2(_05900_),
    .A3(_05902_),
    .B1(_05932_),
    .B2(_05896_),
    .B3(_05891_),
    .ZN(_05933_));
 AOI221_X2 _29396_ (.A(_05929_),
    .B1(_05930_),
    .B2(_05931_),
    .C1(_05716_),
    .C2(_05933_),
    .ZN(_05934_));
 NOR2_X1 _29397_ (.A1(_05927_),
    .A2(_05934_),
    .ZN(_05935_));
 NAND3_X2 _29398_ (.A1(_05862_),
    .A2(_05913_),
    .A3(_05935_),
    .ZN(_05936_));
 XNOR2_X1 _29399_ (.A(_05805_),
    .B(_05936_),
    .ZN(_05937_));
 MUX2_X1 _29400_ (.A(_22406_),
    .B(_05773_),
    .S(_05937_),
    .Z(_05938_));
 MUX2_X1 _29401_ (.A(\g_reduce0[8].adder.x[0] ),
    .B(_05938_),
    .S(_05308_),
    .Z(_05939_));
 OR4_X2 _29402_ (.A1(_05300_),
    .A2(_05301_),
    .A3(_05302_),
    .A4(_05303_),
    .ZN(_05940_));
 CLKBUF_X3 _29403_ (.A(_05940_),
    .Z(_05941_));
 MUX2_X1 _29404_ (.A(\g_reduce0[10].adder.x[0] ),
    .B(_05939_),
    .S(_05941_),
    .Z(_00160_));
 NAND2_X1 _29405_ (.A1(\g_reduce0[10].adder.x[1] ),
    .A2(_05304_),
    .ZN(_05942_));
 NOR4_X4 _29406_ (.A1(\g_reduce0[10].adder.x[11] ),
    .A2(\g_reduce0[10].adder.x[12] ),
    .A3(_05305_),
    .A4(_05306_),
    .ZN(_05943_));
 XNOR2_X1 _29407_ (.A(_22405_),
    .B(_05880_),
    .ZN(_05944_));
 NOR2_X1 _29408_ (.A1(_05943_),
    .A2(_05944_),
    .ZN(_05945_));
 NOR2_X1 _29409_ (.A1(_22406_),
    .A2(_05943_),
    .ZN(_05946_));
 MUX2_X1 _29410_ (.A(_05945_),
    .B(_05946_),
    .S(_05937_),
    .Z(_05947_));
 OAI21_X1 _29411_ (.A(_05941_),
    .B1(_05308_),
    .B2(\g_reduce0[8].adder.x[1] ),
    .ZN(_05948_));
 OAI21_X1 _29412_ (.A(_05942_),
    .B1(_05947_),
    .B2(_05948_),
    .ZN(_00167_));
 NAND2_X1 _29413_ (.A1(\g_reduce0[10].adder.x[2] ),
    .A2(_05304_),
    .ZN(_05949_));
 NOR2_X1 _29414_ (.A1(_05880_),
    .A2(_05912_),
    .ZN(_05950_));
 XNOR2_X1 _29415_ (.A(_05889_),
    .B(_05950_),
    .ZN(_05951_));
 NOR2_X1 _29416_ (.A1(_05943_),
    .A2(_05951_),
    .ZN(_05952_));
 MUX2_X1 _29417_ (.A(_05952_),
    .B(_05945_),
    .S(_05937_),
    .Z(_05953_));
 OAI21_X1 _29418_ (.A(_05941_),
    .B1(_05308_),
    .B2(\g_reduce0[8].adder.x[2] ),
    .ZN(_05954_));
 OAI21_X1 _29419_ (.A(_05949_),
    .B1(_05953_),
    .B2(_05954_),
    .ZN(_00168_));
 NOR2_X2 _29420_ (.A1(_05304_),
    .A2(_05307_),
    .ZN(_05955_));
 AOI22_X1 _29421_ (.A1(\g_reduce0[10].adder.x[3] ),
    .A2(_05304_),
    .B1(_05955_),
    .B2(\g_reduce0[8].adder.x[3] ),
    .ZN(_05956_));
 NOR2_X2 _29422_ (.A1(_05304_),
    .A2(_05943_),
    .ZN(_05957_));
 INV_X1 _29423_ (.A(_05957_),
    .ZN(_05958_));
 NOR2_X1 _29424_ (.A1(_05867_),
    .A2(_05873_),
    .ZN(_05959_));
 INV_X1 _29425_ (.A(_22405_),
    .ZN(_05960_));
 NOR3_X1 _29426_ (.A1(_05960_),
    .A2(_05880_),
    .A3(_05889_),
    .ZN(_05961_));
 XNOR2_X1 _29427_ (.A(_05959_),
    .B(_05961_),
    .ZN(_05962_));
 NOR2_X1 _29428_ (.A1(_05937_),
    .A2(_05962_),
    .ZN(_05963_));
 AOI21_X1 _29429_ (.A(_05963_),
    .B1(_05951_),
    .B2(_05937_),
    .ZN(_05964_));
 OAI21_X1 _29430_ (.A(_05956_),
    .B1(_05958_),
    .B2(_05964_),
    .ZN(_00169_));
 AOI22_X2 _29431_ (.A1(\g_reduce0[10].adder.x[4] ),
    .A2(_05304_),
    .B1(_05955_),
    .B2(\g_reduce0[8].adder.x[4] ),
    .ZN(_05965_));
 OR2_X1 _29432_ (.A1(_05890_),
    .A2(_05912_),
    .ZN(_05966_));
 XNOR2_X1 _29433_ (.A(_05904_),
    .B(_05966_),
    .ZN(_05967_));
 MUX2_X1 _29434_ (.A(_05967_),
    .B(_05962_),
    .S(_05937_),
    .Z(_05968_));
 OAI21_X2 _29435_ (.A(_05965_),
    .B1(_05968_),
    .B2(_05958_),
    .ZN(_00170_));
 NOR2_X1 _29436_ (.A1(\g_reduce0[10].adder.x[5] ),
    .A2(_05941_),
    .ZN(_05969_));
 INV_X1 _29437_ (.A(_05805_),
    .ZN(_05970_));
 OR3_X2 _29438_ (.A1(_05960_),
    .A2(_05890_),
    .A3(_05904_),
    .ZN(_05971_));
 XNOR2_X1 _29439_ (.A(_05827_),
    .B(_05971_),
    .ZN(_05972_));
 OAI221_X1 _29440_ (.A(_05308_),
    .B1(_05970_),
    .B2(_05967_),
    .C1(_05972_),
    .C2(_05937_),
    .ZN(_05973_));
 OAI21_X1 _29441_ (.A(_05973_),
    .B1(_05308_),
    .B2(\g_reduce0[8].adder.x[5] ),
    .ZN(_05974_));
 AOI21_X1 _29442_ (.A(_05969_),
    .B1(_05974_),
    .B2(_05941_),
    .ZN(_00171_));
 NAND2_X1 _29443_ (.A1(\g_reduce0[10].adder.x[6] ),
    .A2(_05304_),
    .ZN(_05975_));
 OAI21_X1 _29444_ (.A(_05941_),
    .B1(_05308_),
    .B2(\g_reduce0[8].adder.x[6] ),
    .ZN(_05976_));
 NOR3_X1 _29445_ (.A1(_05827_),
    .A2(_05904_),
    .A3(_05966_),
    .ZN(_05977_));
 AOI22_X1 _29446_ (.A1(_05801_),
    .A2(_05830_),
    .B1(_05833_),
    .B2(_05746_),
    .ZN(_05978_));
 NAND2_X1 _29447_ (.A1(_05791_),
    .A2(_05931_),
    .ZN(_05979_));
 NAND2_X1 _29448_ (.A1(_05978_),
    .A2(_05979_),
    .ZN(_05980_));
 XNOR2_X1 _29449_ (.A(_05977_),
    .B(_05980_),
    .ZN(_05981_));
 OR2_X1 _29450_ (.A1(_05936_),
    .A2(_05972_),
    .ZN(_05982_));
 AOI21_X1 _29451_ (.A(_05805_),
    .B1(_05981_),
    .B2(_05982_),
    .ZN(_05983_));
 INV_X1 _29452_ (.A(_05936_),
    .ZN(_05984_));
 NOR3_X1 _29453_ (.A1(_05970_),
    .A2(_05984_),
    .A3(_05972_),
    .ZN(_05985_));
 NOR3_X1 _29454_ (.A1(_05943_),
    .A2(_05983_),
    .A3(_05985_),
    .ZN(_05986_));
 OAI21_X1 _29455_ (.A(_05975_),
    .B1(_05976_),
    .B2(_05986_),
    .ZN(_00172_));
 NOR2_X1 _29456_ (.A1(\g_reduce0[10].adder.x[7] ),
    .A2(_05940_),
    .ZN(_05987_));
 NOR2_X1 _29457_ (.A1(_05836_),
    .A2(_05861_),
    .ZN(_05988_));
 OR3_X1 _29458_ (.A1(_05827_),
    .A2(_05834_),
    .A3(_05971_),
    .ZN(_05989_));
 XOR2_X2 _29459_ (.A(_05988_),
    .B(_05989_),
    .Z(_05990_));
 MUX2_X1 _29460_ (.A(_05990_),
    .B(_05981_),
    .S(_05937_),
    .Z(_05991_));
 INV_X1 _29461_ (.A(\g_reduce0[8].adder.x[7] ),
    .ZN(_05992_));
 AOI221_X1 _29462_ (.A(_05987_),
    .B1(_05991_),
    .B2(_05957_),
    .C1(_05955_),
    .C2(_05992_),
    .ZN(_00173_));
 NAND2_X1 _29463_ (.A1(_05862_),
    .A2(_05913_),
    .ZN(_05993_));
 NOR2_X1 _29464_ (.A1(_05934_),
    .A2(_05993_),
    .ZN(_05994_));
 NAND3_X1 _29465_ (.A1(_05994_),
    .A2(_05957_),
    .A3(_05990_),
    .ZN(_05995_));
 NOR2_X1 _29466_ (.A1(_05970_),
    .A2(_05958_),
    .ZN(_05996_));
 OAI21_X1 _29467_ (.A(_05996_),
    .B1(_05990_),
    .B2(_05984_),
    .ZN(_05997_));
 AND2_X1 _29468_ (.A1(_05923_),
    .A2(_05926_),
    .ZN(_05998_));
 OR3_X1 _29469_ (.A1(_05998_),
    .A2(_05917_),
    .A3(_05921_),
    .ZN(_05999_));
 NOR2_X1 _29470_ (.A1(_05999_),
    .A2(_05934_),
    .ZN(_06000_));
 MUX2_X1 _29471_ (.A(_06000_),
    .B(_05934_),
    .S(_05993_),
    .Z(_06001_));
 NAND3_X1 _29472_ (.A1(_05970_),
    .A2(_05957_),
    .A3(_06001_),
    .ZN(_06002_));
 NOR2_X1 _29473_ (.A1(\g_reduce0[10].adder.x[8] ),
    .A2(_05940_),
    .ZN(_06003_));
 INV_X1 _29474_ (.A(\g_reduce0[8].adder.x[8] ),
    .ZN(_06004_));
 AOI21_X1 _29475_ (.A(_06003_),
    .B1(_05955_),
    .B2(_06004_),
    .ZN(_06005_));
 AND4_X1 _29476_ (.A1(_05995_),
    .A2(_05997_),
    .A3(_06002_),
    .A4(_06005_),
    .ZN(_00174_));
 NOR2_X1 _29477_ (.A1(\g_reduce0[10].adder.x[9] ),
    .A2(_05940_),
    .ZN(_06006_));
 NAND3_X1 _29478_ (.A1(_05805_),
    .A2(_05935_),
    .A3(_05971_),
    .ZN(_06007_));
 NAND2_X1 _29479_ (.A1(_05957_),
    .A2(_06007_),
    .ZN(_06008_));
 INV_X1 _29480_ (.A(_05934_),
    .ZN(_06009_));
 XNOR2_X1 _29481_ (.A(_06009_),
    .B(_05993_),
    .ZN(_06010_));
 AOI21_X1 _29482_ (.A(_06008_),
    .B1(_06010_),
    .B2(_05805_),
    .ZN(_06011_));
 NOR2_X1 _29483_ (.A1(_05913_),
    .A2(_05927_),
    .ZN(_06012_));
 AND2_X1 _29484_ (.A1(_05862_),
    .A2(_06009_),
    .ZN(_06013_));
 NOR2_X1 _29485_ (.A1(_05999_),
    .A2(_05971_),
    .ZN(_06014_));
 AOI22_X1 _29486_ (.A1(_05971_),
    .A2(_06012_),
    .B1(_06013_),
    .B2(_06014_),
    .ZN(_06015_));
 OAI21_X1 _29487_ (.A(_06015_),
    .B1(_06013_),
    .B2(_05927_),
    .ZN(_06016_));
 NAND2_X1 _29488_ (.A1(_05970_),
    .A2(_06016_),
    .ZN(_06017_));
 INV_X1 _29489_ (.A(\g_reduce0[8].adder.x[9] ),
    .ZN(_06018_));
 AOI221_X2 _29490_ (.A(_06006_),
    .B1(_06011_),
    .B2(_06017_),
    .C1(_06018_),
    .C2(_05955_),
    .ZN(_00175_));
 INV_X1 _29491_ (.A(_22407_),
    .ZN(_22413_));
 MUX2_X1 _29492_ (.A(\g_reduce0[8].adder.x[10] ),
    .B(_22412_),
    .S(_05308_),
    .Z(_06019_));
 MUX2_X1 _29493_ (.A(\g_reduce0[10].adder.x[10] ),
    .B(_06019_),
    .S(_05941_),
    .Z(_00161_));
 MUX2_X1 _29494_ (.A(_05300_),
    .B(_22420_),
    .S(_05308_),
    .Z(_06020_));
 MUX2_X1 _29495_ (.A(\g_reduce0[10].adder.x[11] ),
    .B(_06020_),
    .S(_05941_),
    .Z(_00162_));
 XOR2_X1 _29496_ (.A(_14192_),
    .B(_22424_),
    .Z(_06021_));
 MUX2_X2 _29497_ (.A(_22285_),
    .B(_00598_),
    .S(_05367_),
    .Z(_06022_));
 NAND2_X1 _29498_ (.A1(_05714_),
    .A2(_22414_),
    .ZN(_06023_));
 XOR2_X1 _29499_ (.A(_06022_),
    .B(_06023_),
    .Z(_06024_));
 MUX2_X1 _29500_ (.A(_06021_),
    .B(_06024_),
    .S(_05746_),
    .Z(_06025_));
 XOR2_X1 _29501_ (.A(_22419_),
    .B(_06025_),
    .Z(_06026_));
 MUX2_X1 _29502_ (.A(_05301_),
    .B(_06026_),
    .S(_05307_),
    .Z(_06027_));
 MUX2_X1 _29503_ (.A(\g_reduce0[10].adder.x[12] ),
    .B(_06027_),
    .S(_05941_),
    .Z(_00163_));
 INV_X1 _29504_ (.A(_14194_),
    .ZN(_14191_));
 INV_X1 _29505_ (.A(_22416_),
    .ZN(_06028_));
 INV_X1 _29506_ (.A(_22417_),
    .ZN(_06029_));
 OAI21_X1 _29507_ (.A(_06028_),
    .B1(_06029_),
    .B2(_14194_),
    .ZN(_06030_));
 AOI21_X1 _29508_ (.A(_22423_),
    .B1(_06030_),
    .B2(_22424_),
    .ZN(_06031_));
 XNOR2_X1 _29509_ (.A(_22428_),
    .B(_06031_),
    .ZN(_06032_));
 MUX2_X2 _29510_ (.A(_22282_),
    .B(_00601_),
    .S(_05367_),
    .Z(_06033_));
 MUX2_X1 _29511_ (.A(_22288_),
    .B(_00593_),
    .S(_05367_),
    .Z(_06034_));
 NOR4_X1 _29512_ (.A1(_05733_),
    .A2(_22407_),
    .A3(_06022_),
    .A4(_06034_),
    .ZN(_06035_));
 XNOR2_X1 _29513_ (.A(_06033_),
    .B(_06035_),
    .ZN(_06036_));
 MUX2_X1 _29514_ (.A(_06032_),
    .B(_06036_),
    .S(_05746_),
    .Z(_06037_));
 NAND2_X1 _29515_ (.A1(_05714_),
    .A2(_22415_),
    .ZN(_06038_));
 OAI21_X1 _29516_ (.A(_06038_),
    .B1(_06034_),
    .B2(_05714_),
    .ZN(_06039_));
 MUX2_X1 _29517_ (.A(_14193_),
    .B(_06039_),
    .S(_05746_),
    .Z(_22418_));
 NAND3_X1 _29518_ (.A1(_22411_),
    .A2(_06025_),
    .A3(_22418_),
    .ZN(_06040_));
 XNOR2_X1 _29519_ (.A(_06037_),
    .B(_06040_),
    .ZN(_06041_));
 MUX2_X1 _29520_ (.A(\g_reduce0[8].adder.x[13] ),
    .B(_06041_),
    .S(_05307_),
    .Z(_06042_));
 MUX2_X1 _29521_ (.A(\g_reduce0[10].adder.x[13] ),
    .B(_06042_),
    .S(_05941_),
    .Z(_00164_));
 NOR4_X2 _29522_ (.A1(_05716_),
    .A2(_06022_),
    .A3(_06023_),
    .A4(_06033_),
    .ZN(_06043_));
 AOI21_X1 _29523_ (.A(_22423_),
    .B1(_22424_),
    .B2(_14192_),
    .ZN(_06044_));
 INV_X1 _29524_ (.A(_06044_),
    .ZN(_06045_));
 AOI21_X1 _29525_ (.A(_22427_),
    .B1(_06045_),
    .B2(_22428_),
    .ZN(_06046_));
 AOI21_X2 _29526_ (.A(_06043_),
    .B1(_06046_),
    .B2(_05716_),
    .ZN(_06047_));
 NAND3_X1 _29527_ (.A1(_22419_),
    .A2(_06025_),
    .A3(_06037_),
    .ZN(_06048_));
 XOR2_X2 _29528_ (.A(_06047_),
    .B(_06048_),
    .Z(_06049_));
 OAI21_X1 _29529_ (.A(_05308_),
    .B1(_05354_),
    .B2(_06049_),
    .ZN(_06050_));
 OAI21_X1 _29530_ (.A(_05940_),
    .B1(_05319_),
    .B2(_06049_),
    .ZN(_06051_));
 MUX2_X1 _29531_ (.A(_05302_),
    .B(_05305_),
    .S(_05354_),
    .Z(_06052_));
 OAI21_X1 _29532_ (.A(_05307_),
    .B1(_05940_),
    .B2(_05305_),
    .ZN(_06053_));
 INV_X1 _29533_ (.A(_05302_),
    .ZN(_06054_));
 AOI21_X1 _29534_ (.A(_06052_),
    .B1(_06053_),
    .B2(_06054_),
    .ZN(_06055_));
 AOI222_X2 _29535_ (.A1(_05302_),
    .A2(_06050_),
    .B1(_06051_),
    .B2(_05305_),
    .C1(_06049_),
    .C2(_06055_),
    .ZN(_06056_));
 INV_X1 _29536_ (.A(_06056_),
    .ZN(_00165_));
 CLKBUF_X2 _29537_ (.A(\g_reduce0[12].adder.x[11] ),
    .Z(_06057_));
 CLKBUF_X2 _29538_ (.A(\g_reduce0[12].adder.x[12] ),
    .Z(_06058_));
 BUF_X2 _29539_ (.A(\g_reduce0[12].adder.x[14] ),
    .Z(_06059_));
 OR2_X1 _29540_ (.A1(\g_reduce0[12].adder.x[10] ),
    .A2(\g_reduce0[12].adder.x[13] ),
    .ZN(_06060_));
 OR4_X2 _29541_ (.A1(_06057_),
    .A2(_06058_),
    .A3(_06059_),
    .A4(_06060_),
    .ZN(_06061_));
 BUF_X2 _29542_ (.A(\g_reduce0[14].adder.x[14] ),
    .Z(_06062_));
 OR2_X2 _29543_ (.A1(\g_reduce0[14].adder.x[10] ),
    .A2(\g_reduce0[14].adder.x[13] ),
    .ZN(_06063_));
 NOR4_X4 _29544_ (.A1(\g_reduce0[14].adder.x[11] ),
    .A2(\g_reduce0[14].adder.x[12] ),
    .A3(_06062_),
    .A4(_06063_),
    .ZN(_06064_));
 OR2_X1 _29545_ (.A1(_22475_),
    .A2(_22430_),
    .ZN(_06065_));
 INV_X1 _29546_ (.A(_22436_),
    .ZN(_06066_));
 INV_X1 _29547_ (.A(_22437_),
    .ZN(_06067_));
 OAI21_X1 _29548_ (.A(_06066_),
    .B1(_22469_),
    .B2(_06067_),
    .ZN(_06068_));
 BUF_X4 _29549_ (.A(_22431_),
    .Z(_06069_));
 BUF_X4 _29550_ (.A(_22434_),
    .Z(_06070_));
 AND2_X1 _29551_ (.A1(_06069_),
    .A2(_06070_),
    .ZN(_06071_));
 AOI221_X4 _29552_ (.A(_06065_),
    .B1(_06068_),
    .B2(_06071_),
    .C1(_06069_),
    .C2(_22433_),
    .ZN(_06072_));
 INV_X2 _29553_ (.A(_22476_),
    .ZN(_06073_));
 CLKBUF_X3 _29554_ (.A(_22470_),
    .Z(_06074_));
 INV_X2 _29555_ (.A(_06074_),
    .ZN(_06075_));
 NAND2_X1 _29556_ (.A1(_06069_),
    .A2(_06070_),
    .ZN(_06076_));
 NOR4_X1 _29557_ (.A1(_06073_),
    .A2(_06075_),
    .A3(_06067_),
    .A4(_06076_),
    .ZN(_06077_));
 NOR2_X1 _29558_ (.A1(_22476_),
    .A2(_22475_),
    .ZN(_06078_));
 OR2_X2 _29559_ (.A1(_06077_),
    .A2(_06078_),
    .ZN(_06079_));
 AOI21_X1 _29560_ (.A(_22439_),
    .B1(_22442_),
    .B2(_22440_),
    .ZN(_06080_));
 NAND2_X1 _29561_ (.A1(_22440_),
    .A2(_22443_),
    .ZN(_06081_));
 AOI21_X1 _29562_ (.A(_22445_),
    .B1(_22446_),
    .B2(_22448_),
    .ZN(_06082_));
 OAI21_X1 _29563_ (.A(_06080_),
    .B1(_06081_),
    .B2(_06082_),
    .ZN(_06083_));
 AND4_X1 _29564_ (.A1(_22440_),
    .A2(_22443_),
    .A3(_22446_),
    .A4(_22449_),
    .ZN(_06084_));
 AND3_X1 _29565_ (.A1(_22452_),
    .A2(_22455_),
    .A3(_22458_),
    .ZN(_06085_));
 AND3_X1 _29566_ (.A1(_22461_),
    .A2(_06084_),
    .A3(_06085_),
    .ZN(_06086_));
 INV_X1 _29567_ (.A(_22463_),
    .ZN(_06087_));
 INV_X1 _29568_ (.A(_22464_),
    .ZN(_06088_));
 OAI21_X1 _29569_ (.A(_06087_),
    .B1(_22466_),
    .B2(_06088_),
    .ZN(_06089_));
 INV_X1 _29570_ (.A(_22451_),
    .ZN(_06090_));
 NAND3_X1 _29571_ (.A1(_22452_),
    .A2(_22455_),
    .A3(_22458_),
    .ZN(_06091_));
 INV_X1 _29572_ (.A(_22460_),
    .ZN(_06092_));
 AOI21_X1 _29573_ (.A(_22454_),
    .B1(_22457_),
    .B2(_22455_),
    .ZN(_06093_));
 INV_X1 _29574_ (.A(_22452_),
    .ZN(_06094_));
 OAI221_X2 _29575_ (.A(_06090_),
    .B1(_06091_),
    .B2(_06092_),
    .C1(_06093_),
    .C2(_06094_),
    .ZN(_06095_));
 AOI221_X2 _29576_ (.A(_06083_),
    .B1(_06086_),
    .B2(_06089_),
    .C1(_06095_),
    .C2(_06084_),
    .ZN(_06096_));
 NAND3_X1 _29577_ (.A1(_22461_),
    .A2(_06084_),
    .A3(_06085_),
    .ZN(_06097_));
 NAND2_X1 _29578_ (.A1(_22464_),
    .A2(_22467_),
    .ZN(_06098_));
 OAI21_X1 _29579_ (.A(_06077_),
    .B1(_06097_),
    .B2(_06098_),
    .ZN(_06099_));
 OAI22_X4 _29580_ (.A1(_06072_),
    .A2(_06079_),
    .B1(_06096_),
    .B2(_06099_),
    .ZN(_06100_));
 CLKBUF_X3 _29581_ (.A(_06100_),
    .Z(_06101_));
 CLKBUF_X3 _29582_ (.A(_06101_),
    .Z(_06102_));
 OAI21_X1 _29583_ (.A(_06061_),
    .B1(_06064_),
    .B2(_06102_),
    .ZN(_06103_));
 MUX2_X1 _29584_ (.A(\g_reduce0[12].adder.x[15] ),
    .B(\g_reduce0[14].adder.x[15] ),
    .S(_06103_),
    .Z(_00182_));
 INV_X1 _29585_ (.A(_00604_),
    .ZN(_06104_));
 INV_X1 _29586_ (.A(_22468_),
    .ZN(_06105_));
 MUX2_X2 _29587_ (.A(_06104_),
    .B(_06105_),
    .S(_06102_),
    .Z(_19424_));
 INV_X1 _29588_ (.A(_19424_),
    .ZN(_22554_));
 MUX2_X2 _29589_ (.A(_22435_),
    .B(_00607_),
    .S(_06102_),
    .Z(_14205_));
 NOR2_X1 _29590_ (.A1(\g_reduce0[12].adder.x[13] ),
    .A2(_22429_),
    .ZN(_06106_));
 NOR2_X1 _29591_ (.A1(\g_reduce0[14].adder.x[13] ),
    .A2(_00615_),
    .ZN(_06107_));
 MUX2_X1 _29592_ (.A(_06106_),
    .B(_06107_),
    .S(_06100_),
    .Z(_06108_));
 NOR2_X1 _29593_ (.A1(_06058_),
    .A2(_22432_),
    .ZN(_06109_));
 NOR2_X1 _29594_ (.A1(\g_reduce0[14].adder.x[12] ),
    .A2(_00612_),
    .ZN(_06110_));
 MUX2_X2 _29595_ (.A(_06109_),
    .B(_06110_),
    .S(_06100_),
    .Z(_06111_));
 NOR2_X1 _29596_ (.A1(_06057_),
    .A2(_22435_),
    .ZN(_06112_));
 OR2_X1 _29597_ (.A1(_22472_),
    .A2(_06112_),
    .ZN(_06113_));
 NOR2_X1 _29598_ (.A1(\g_reduce0[14].adder.x[11] ),
    .A2(_00607_),
    .ZN(_06114_));
 OR2_X1 _29599_ (.A1(_22472_),
    .A2(_06114_),
    .ZN(_06115_));
 MUX2_X2 _29600_ (.A(_06113_),
    .B(_06115_),
    .S(_06100_),
    .Z(_06116_));
 OR4_X2 _29601_ (.A1(_22476_),
    .A2(_06108_),
    .A3(_06111_),
    .A4(_06116_),
    .ZN(_06117_));
 INV_X1 _29602_ (.A(_06069_),
    .ZN(_06118_));
 NOR2_X2 _29603_ (.A1(_06073_),
    .A2(_06118_),
    .ZN(_06119_));
 AND2_X1 _29604_ (.A1(_06070_),
    .A2(_06119_),
    .ZN(_06120_));
 AOI22_X4 _29605_ (.A1(_06111_),
    .A2(_06119_),
    .B1(_06120_),
    .B2(_06116_),
    .ZN(_06121_));
 OR4_X2 _29606_ (.A1(_22476_),
    .A2(_06070_),
    .A3(_06108_),
    .A4(_06111_),
    .ZN(_06122_));
 NAND2_X1 _29607_ (.A1(_06073_),
    .A2(_06118_),
    .ZN(_06123_));
 MUX2_X1 _29608_ (.A(_06123_),
    .B(_06073_),
    .S(_06108_),
    .Z(_06124_));
 NAND4_X4 _29609_ (.A1(_06117_),
    .A2(_06121_),
    .A3(_06122_),
    .A4(_06124_),
    .ZN(_06125_));
 XOR2_X2 _29610_ (.A(_06070_),
    .B(_06116_),
    .Z(_06126_));
 CLKBUF_X3 _29611_ (.A(_06075_),
    .Z(_06127_));
 MUX2_X1 _29612_ (.A(_00614_),
    .B(_22441_),
    .S(_06101_),
    .Z(_06128_));
 MUX2_X1 _29613_ (.A(_00613_),
    .B(_22438_),
    .S(_06101_),
    .Z(_06129_));
 MUX2_X1 _29614_ (.A(_06128_),
    .B(_06129_),
    .S(_06127_),
    .Z(_06130_));
 CLKBUF_X3 _29615_ (.A(_22473_),
    .Z(_06131_));
 INV_X2 _29616_ (.A(_06131_),
    .ZN(_06132_));
 MUX2_X1 _29617_ (.A(_06127_),
    .B(_06130_),
    .S(_06132_),
    .Z(_06133_));
 MUX2_X1 _29618_ (.A(_22465_),
    .B(_00603_),
    .S(_06101_),
    .Z(_06134_));
 MUX2_X1 _29619_ (.A(_00606_),
    .B(_22459_),
    .S(_06100_),
    .Z(_06135_));
 MUX2_X1 _29620_ (.A(_06134_),
    .B(_06135_),
    .S(_06131_),
    .Z(_06136_));
 MUX2_X1 _29621_ (.A(_00602_),
    .B(_22462_),
    .S(_06102_),
    .Z(_06137_));
 MUX2_X1 _29622_ (.A(_00605_),
    .B(_22456_),
    .S(_06102_),
    .Z(_06138_));
 MUX2_X1 _29623_ (.A(_06137_),
    .B(_06138_),
    .S(_06131_),
    .Z(_06139_));
 MUX2_X1 _29624_ (.A(_06136_),
    .B(_06139_),
    .S(_06127_),
    .Z(_06140_));
 MUX2_X2 _29625_ (.A(_06112_),
    .B(_06114_),
    .S(_06100_),
    .Z(_06141_));
 NOR2_X1 _29626_ (.A1(_06104_),
    .A2(_22468_),
    .ZN(_06142_));
 OAI211_X2 _29627_ (.A(_06099_),
    .B(_06142_),
    .C1(_06072_),
    .C2(_06079_),
    .ZN(_06143_));
 OR4_X1 _29628_ (.A1(_00604_),
    .A2(_06105_),
    .A3(_06096_),
    .A4(_06099_),
    .ZN(_06144_));
 OAI211_X2 _29629_ (.A(_06096_),
    .B(_06142_),
    .C1(_06072_),
    .C2(_06079_),
    .ZN(_06145_));
 OR4_X1 _29630_ (.A1(_00604_),
    .A2(_06105_),
    .A3(_06072_),
    .A4(_06079_),
    .ZN(_06146_));
 AND4_X2 _29631_ (.A1(_06143_),
    .A2(_06144_),
    .A3(_06145_),
    .A4(_06146_),
    .ZN(_22471_));
 OR4_X2 _29632_ (.A1(_06069_),
    .A2(_06111_),
    .A3(_06141_),
    .A4(_22471_),
    .ZN(_06147_));
 NOR2_X1 _29633_ (.A1(_06067_),
    .A2(_06076_),
    .ZN(_06148_));
 AOI22_X4 _29634_ (.A1(_06071_),
    .A2(_06141_),
    .B1(_22471_),
    .B2(_06148_),
    .ZN(_06149_));
 OR4_X2 _29635_ (.A1(_06069_),
    .A2(_22437_),
    .A3(_06111_),
    .A4(_06141_),
    .ZN(_06150_));
 OR2_X1 _29636_ (.A1(_06069_),
    .A2(_06070_),
    .ZN(_06151_));
 MUX2_X1 _29637_ (.A(_06151_),
    .B(_06118_),
    .S(_06111_),
    .Z(_06152_));
 NAND4_X4 _29638_ (.A1(_06147_),
    .A2(_06149_),
    .A3(_06150_),
    .A4(_06152_),
    .ZN(_06153_));
 MUX2_X1 _29639_ (.A(_06133_),
    .B(_06140_),
    .S(_06153_),
    .Z(_06154_));
 MUX2_X1 _29640_ (.A(_00611_),
    .B(_22447_),
    .S(_06101_),
    .Z(_06155_));
 MUX2_X1 _29641_ (.A(_00610_),
    .B(_22444_),
    .S(_06101_),
    .Z(_06156_));
 MUX2_X1 _29642_ (.A(_06155_),
    .B(_06156_),
    .S(_06127_),
    .Z(_06157_));
 MUX2_X1 _29643_ (.A(_00609_),
    .B(_22453_),
    .S(_06101_),
    .Z(_06158_));
 MUX2_X1 _29644_ (.A(_00608_),
    .B(_22450_),
    .S(_06102_),
    .Z(_06159_));
 MUX2_X1 _29645_ (.A(_06158_),
    .B(_06159_),
    .S(_06127_),
    .Z(_06160_));
 MUX2_X1 _29646_ (.A(_06157_),
    .B(_06160_),
    .S(_06132_),
    .Z(_06161_));
 NAND2_X1 _29647_ (.A1(_06126_),
    .A2(_06153_),
    .ZN(_06162_));
 OAI22_X1 _29648_ (.A1(_06126_),
    .A2(_06154_),
    .B1(_06161_),
    .B2(_06162_),
    .ZN(_06163_));
 NAND2_X1 _29649_ (.A1(_06125_),
    .A2(_06163_),
    .ZN(_22540_));
 INV_X1 _29650_ (.A(_22540_),
    .ZN(_22538_));
 AND4_X1 _29651_ (.A1(_06117_),
    .A2(_06121_),
    .A3(_06122_),
    .A4(_06124_),
    .ZN(_06164_));
 BUF_X4 _29652_ (.A(_06164_),
    .Z(_06165_));
 MUX2_X1 _29653_ (.A(_06128_),
    .B(_06155_),
    .S(_06132_),
    .Z(_06166_));
 MUX2_X1 _29654_ (.A(_06156_),
    .B(_06159_),
    .S(_06132_),
    .Z(_06167_));
 MUX2_X1 _29655_ (.A(_06166_),
    .B(_06167_),
    .S(_06074_),
    .Z(_06168_));
 NOR2_X1 _29656_ (.A1(_06162_),
    .A2(_06168_),
    .ZN(_06169_));
 AND4_X1 _29657_ (.A1(_06147_),
    .A2(_06149_),
    .A3(_06150_),
    .A4(_06152_),
    .ZN(_06170_));
 BUF_X4 _29658_ (.A(_06170_),
    .Z(_06171_));
 AOI21_X2 _29659_ (.A(_06131_),
    .B1(_06129_),
    .B2(_06074_),
    .ZN(_06172_));
 NAND2_X1 _29660_ (.A1(_06171_),
    .A2(_06172_),
    .ZN(_06173_));
 MUX2_X1 _29661_ (.A(_06135_),
    .B(_06158_),
    .S(_06131_),
    .Z(_06174_));
 MUX2_X1 _29662_ (.A(_06139_),
    .B(_06174_),
    .S(_06127_),
    .Z(_06175_));
 OAI21_X1 _29663_ (.A(_06173_),
    .B1(_06175_),
    .B2(_06171_),
    .ZN(_06176_));
 XNOR2_X1 _29664_ (.A(_06070_),
    .B(_06116_),
    .ZN(_06177_));
 BUF_X4 _29665_ (.A(_06177_),
    .Z(_06178_));
 AOI21_X1 _29666_ (.A(_06169_),
    .B1(_06176_),
    .B2(_06178_),
    .ZN(_06179_));
 OR2_X1 _29667_ (.A1(_06165_),
    .A2(_06179_),
    .ZN(_14201_));
 INV_X1 _29668_ (.A(_14201_),
    .ZN(_14197_));
 NOR2_X2 _29669_ (.A1(_06165_),
    .A2(_06171_),
    .ZN(_06180_));
 NAND3_X2 _29670_ (.A1(_06178_),
    .A2(_06172_),
    .A3(_06180_),
    .ZN(_22492_));
 INV_X1 _29671_ (.A(_22492_),
    .ZN(_22496_));
 NAND2_X1 _29672_ (.A1(_06125_),
    .A2(_06153_),
    .ZN(_06181_));
 OR3_X1 _29673_ (.A1(_06126_),
    .A2(_06133_),
    .A3(_06181_),
    .ZN(_22486_));
 INV_X1 _29674_ (.A(_22486_),
    .ZN(_22489_));
 NOR2_X1 _29675_ (.A1(_06074_),
    .A2(_06131_),
    .ZN(_06182_));
 NOR2_X1 _29676_ (.A1(_06075_),
    .A2(_06132_),
    .ZN(_06183_));
 AOI22_X2 _29677_ (.A1(_06128_),
    .A2(_06182_),
    .B1(_06183_),
    .B2(_06129_),
    .ZN(_06184_));
 NOR2_X2 _29678_ (.A1(_06075_),
    .A2(_06131_),
    .ZN(_06185_));
 NAND2_X1 _29679_ (.A1(_06156_),
    .A2(_06185_),
    .ZN(_06186_));
 AND2_X1 _29680_ (.A1(_06184_),
    .A2(_06186_),
    .ZN(_06187_));
 NAND3_X1 _29681_ (.A1(_06178_),
    .A2(_06180_),
    .A3(_06187_),
    .ZN(_22520_));
 INV_X1 _29682_ (.A(_22520_),
    .ZN(_22524_));
 NAND2_X1 _29683_ (.A1(_06126_),
    .A2(_06185_),
    .ZN(_06188_));
 MUX2_X1 _29684_ (.A(_06130_),
    .B(_06157_),
    .S(_06132_),
    .Z(_06189_));
 OAI21_X1 _29685_ (.A(_06188_),
    .B1(_06189_),
    .B2(_06126_),
    .ZN(_06190_));
 NAND2_X1 _29686_ (.A1(_06180_),
    .A2(_06190_),
    .ZN(_22499_));
 INV_X1 _29687_ (.A(_22499_),
    .ZN(_22503_));
 NAND2_X1 _29688_ (.A1(_06126_),
    .A2(_06172_),
    .ZN(_06191_));
 OAI21_X1 _29689_ (.A(_06191_),
    .B1(_06168_),
    .B2(_06126_),
    .ZN(_06192_));
 AND2_X1 _29690_ (.A1(_06180_),
    .A2(_06192_),
    .ZN(_22507_));
 INV_X1 _29691_ (.A(_22507_),
    .ZN(_22510_));
 MUX2_X1 _29692_ (.A(_06133_),
    .B(_06161_),
    .S(_06178_),
    .Z(_06193_));
 NOR2_X1 _29693_ (.A1(_06181_),
    .A2(_06193_),
    .ZN(_22513_));
 INV_X1 _29694_ (.A(_22513_),
    .ZN(_22517_));
 INV_X1 _29695_ (.A(_06182_),
    .ZN(_06194_));
 MUX2_X1 _29696_ (.A(_00605_),
    .B(_00608_),
    .S(_22473_),
    .Z(_06195_));
 MUX2_X1 _29697_ (.A(_22456_),
    .B(_22450_),
    .S(_22473_),
    .Z(_06196_));
 MUX2_X1 _29698_ (.A(_06195_),
    .B(_06196_),
    .S(_06101_),
    .Z(_06197_));
 OAI22_X2 _29699_ (.A1(_06158_),
    .A2(_06194_),
    .B1(_06197_),
    .B2(_06127_),
    .ZN(_06198_));
 NOR3_X2 _29700_ (.A1(_06074_),
    .A2(_06132_),
    .A3(_06155_),
    .ZN(_06199_));
 OAI21_X1 _29701_ (.A(_06178_),
    .B1(_06198_),
    .B2(_06199_),
    .ZN(_06200_));
 NAND2_X1 _29702_ (.A1(_06126_),
    .A2(_06187_),
    .ZN(_06201_));
 NAND2_X1 _29703_ (.A1(_06200_),
    .A2(_06201_),
    .ZN(_06202_));
 AND2_X1 _29704_ (.A1(_06180_),
    .A2(_06202_),
    .ZN(_22531_));
 INV_X1 _29705_ (.A(_22531_),
    .ZN(_22534_));
 NOR2_X1 _29706_ (.A1(_06162_),
    .A2(_06189_),
    .ZN(_06203_));
 OR3_X1 _29707_ (.A1(_06074_),
    .A2(_06171_),
    .A3(_06197_),
    .ZN(_06204_));
 MUX2_X1 _29708_ (.A(_06131_),
    .B(_06174_),
    .S(_06153_),
    .Z(_06205_));
 OAI21_X1 _29709_ (.A(_06204_),
    .B1(_06205_),
    .B2(_06127_),
    .ZN(_06206_));
 AOI21_X1 _29710_ (.A(_06203_),
    .B1(_06206_),
    .B2(_06178_),
    .ZN(_06207_));
 OR2_X1 _29711_ (.A1(_06165_),
    .A2(_06207_),
    .ZN(_22527_));
 INV_X1 _29712_ (.A(_22527_),
    .ZN(_22481_));
 XNOR2_X2 _29713_ (.A(\g_reduce0[14].adder.x[15] ),
    .B(\g_reduce0[12].adder.x[15] ),
    .ZN(_06208_));
 BUF_X4 _29714_ (.A(_06208_),
    .Z(_06209_));
 BUF_X4 _29715_ (.A(_06209_),
    .Z(_06210_));
 BUF_X2 _29716_ (.A(_22495_),
    .Z(_06211_));
 BUF_X1 _29717_ (.A(_22488_),
    .Z(_06212_));
 INV_X1 _29718_ (.A(_06212_),
    .ZN(_06213_));
 CLKBUF_X3 _29719_ (.A(_22502_),
    .Z(_06214_));
 BUF_X2 _29720_ (.A(_22523_),
    .Z(_06215_));
 BUF_X2 _29721_ (.A(_22509_),
    .Z(_06216_));
 INV_X1 _29722_ (.A(_06216_),
    .ZN(_06217_));
 BUF_X2 _29723_ (.A(_22516_),
    .Z(_06218_));
 NOR2_X1 _29724_ (.A1(_06218_),
    .A2(_22515_),
    .ZN(_06219_));
 NOR2_X1 _29725_ (.A1(_06217_),
    .A2(_06219_),
    .ZN(_06220_));
 NOR2_X1 _29726_ (.A1(_22508_),
    .A2(_06220_),
    .ZN(_06221_));
 OR3_X1 _29727_ (.A1(_22508_),
    .A2(_22515_),
    .A3(_22532_),
    .ZN(_06222_));
 INV_X1 _29728_ (.A(_22483_),
    .ZN(_06223_));
 INV_X1 _29729_ (.A(_22484_),
    .ZN(_06224_));
 AOI21_X1 _29730_ (.A(_22477_),
    .B1(_14195_),
    .B2(_22478_),
    .ZN(_06225_));
 OAI21_X2 _29731_ (.A(_06223_),
    .B1(_06224_),
    .B2(_06225_),
    .ZN(_06226_));
 BUF_X2 _29732_ (.A(_22533_),
    .Z(_06227_));
 AOI21_X2 _29733_ (.A(_06222_),
    .B1(_06226_),
    .B2(_06227_),
    .ZN(_06228_));
 NOR4_X2 _29734_ (.A1(_06214_),
    .A2(_06215_),
    .A3(_06221_),
    .A4(_06228_),
    .ZN(_06229_));
 INV_X1 _29735_ (.A(_22525_),
    .ZN(_06230_));
 INV_X1 _29736_ (.A(_22504_),
    .ZN(_06231_));
 OAI21_X1 _29737_ (.A(_06230_),
    .B1(_06231_),
    .B2(_06215_),
    .ZN(_06232_));
 OAI21_X1 _29738_ (.A(_06213_),
    .B1(_06229_),
    .B2(_06232_),
    .ZN(_06233_));
 INV_X1 _29739_ (.A(_22490_),
    .ZN(_06234_));
 AOI21_X2 _29740_ (.A(_06211_),
    .B1(_06233_),
    .B2(_06234_),
    .ZN(_06235_));
 OAI21_X4 _29741_ (.A(_06210_),
    .B1(_06235_),
    .B2(_22497_),
    .ZN(_06236_));
 AOI21_X1 _29742_ (.A(_22522_),
    .B1(_22501_),
    .B2(_06215_),
    .ZN(_06237_));
 INV_X1 _29743_ (.A(_22518_),
    .ZN(_06238_));
 AOI21_X1 _29744_ (.A(_06216_),
    .B1(_06218_),
    .B2(_06238_),
    .ZN(_06239_));
 NOR2_X1 _29745_ (.A1(_22511_),
    .A2(_06239_),
    .ZN(_06240_));
 INV_X1 _29746_ (.A(_22511_),
    .ZN(_06241_));
 INV_X1 _29747_ (.A(_22535_),
    .ZN(_06242_));
 NAND3_X1 _29748_ (.A1(_06241_),
    .A2(_06238_),
    .A3(_06242_),
    .ZN(_06243_));
 INV_X1 _29749_ (.A(_22528_),
    .ZN(_06244_));
 INV_X1 _29750_ (.A(_22529_),
    .ZN(_06245_));
 AOI21_X1 _29751_ (.A(_22479_),
    .B1(_14200_),
    .B2(_22480_),
    .ZN(_06246_));
 OAI21_X2 _29752_ (.A(_06244_),
    .B1(_06245_),
    .B2(_06246_),
    .ZN(_06247_));
 INV_X1 _29753_ (.A(_06227_),
    .ZN(_06248_));
 AOI21_X1 _29754_ (.A(_06243_),
    .B1(_06247_),
    .B2(_06248_),
    .ZN(_06249_));
 NAND2_X1 _29755_ (.A1(_06214_),
    .A2(_06215_),
    .ZN(_06250_));
 OR3_X1 _29756_ (.A1(_06240_),
    .A2(_06249_),
    .A3(_06250_),
    .ZN(_06251_));
 AOI21_X1 _29757_ (.A(_06213_),
    .B1(_06237_),
    .B2(_06251_),
    .ZN(_06252_));
 OAI21_X1 _29758_ (.A(_06211_),
    .B1(_22487_),
    .B2(_06252_),
    .ZN(_06253_));
 INV_X1 _29759_ (.A(_22494_),
    .ZN(_06254_));
 AOI21_X1 _29760_ (.A(_06210_),
    .B1(_06253_),
    .B2(_06254_),
    .ZN(_06255_));
 NAND2_X2 _29761_ (.A1(_06178_),
    .A2(_06185_),
    .ZN(_06256_));
 OR4_X2 _29762_ (.A1(_06165_),
    .A2(_06171_),
    .A3(_06255_),
    .A4(_06256_),
    .ZN(_06257_));
 NAND2_X2 _29763_ (.A1(_06236_),
    .A2(_06257_),
    .ZN(_06258_));
 AOI21_X1 _29764_ (.A(_06215_),
    .B1(_06231_),
    .B2(_06214_),
    .ZN(_06259_));
 OR2_X2 _29765_ (.A1(_22525_),
    .A2(_06259_),
    .ZN(_06260_));
 NOR3_X1 _29766_ (.A1(_22525_),
    .A2(_22504_),
    .A3(_22508_),
    .ZN(_06261_));
 INV_X1 _29767_ (.A(_22532_),
    .ZN(_06262_));
 AOI21_X1 _29768_ (.A(_22483_),
    .B1(_14198_),
    .B2(_22484_),
    .ZN(_06263_));
 OAI21_X2 _29769_ (.A(_06262_),
    .B1(_06263_),
    .B2(_06248_),
    .ZN(_06264_));
 AOI21_X1 _29770_ (.A(_22515_),
    .B1(_06264_),
    .B2(_06218_),
    .ZN(_06265_));
 OAI21_X2 _29771_ (.A(_06261_),
    .B1(_06265_),
    .B2(_06217_),
    .ZN(_06266_));
 AND4_X2 _29772_ (.A1(_06212_),
    .A2(_06209_),
    .A3(_06260_),
    .A4(_06266_),
    .ZN(_06267_));
 NAND2_X1 _29773_ (.A1(_06213_),
    .A2(_06209_),
    .ZN(_06268_));
 AOI21_X4 _29774_ (.A(_06268_),
    .B1(_06266_),
    .B2(_06260_),
    .ZN(_06269_));
 XOR2_X2 _29775_ (.A(\g_reduce0[14].adder.x[15] ),
    .B(\g_reduce0[12].adder.x[15] ),
    .Z(_06270_));
 BUF_X4 _29776_ (.A(_06270_),
    .Z(_06271_));
 NAND2_X1 _29777_ (.A1(_06212_),
    .A2(_06271_),
    .ZN(_06272_));
 AND2_X1 _29778_ (.A1(_06241_),
    .A2(_06237_),
    .ZN(_06273_));
 AOI21_X1 _29779_ (.A(_22528_),
    .B1(_14202_),
    .B2(_22529_),
    .ZN(_06274_));
 OAI21_X1 _29780_ (.A(_06242_),
    .B1(_06274_),
    .B2(_06227_),
    .ZN(_06275_));
 INV_X1 _29781_ (.A(_06218_),
    .ZN(_06276_));
 AOI21_X2 _29782_ (.A(_22518_),
    .B1(_06275_),
    .B2(_06276_),
    .ZN(_06277_));
 OAI21_X2 _29783_ (.A(_06273_),
    .B1(_06277_),
    .B2(_06216_),
    .ZN(_06278_));
 INV_X1 _29784_ (.A(_22522_),
    .ZN(_06279_));
 OAI21_X1 _29785_ (.A(_06215_),
    .B1(_22501_),
    .B2(_06214_),
    .ZN(_06280_));
 NAND2_X2 _29786_ (.A1(_06279_),
    .A2(_06280_),
    .ZN(_06281_));
 AOI21_X4 _29787_ (.A(_06272_),
    .B1(_06278_),
    .B2(_06281_),
    .ZN(_06282_));
 AND4_X2 _29788_ (.A1(_06213_),
    .A2(_06271_),
    .A3(_06281_),
    .A4(_06278_),
    .ZN(_06283_));
 NOR4_X4 _29789_ (.A1(_06267_),
    .A2(_06269_),
    .A3(_06282_),
    .A4(_06283_),
    .ZN(_06284_));
 BUF_X4 _29790_ (.A(_06284_),
    .Z(_06285_));
 OAI21_X2 _29791_ (.A(_06241_),
    .B1(_06216_),
    .B2(_06277_),
    .ZN(_06286_));
 OR2_X1 _29792_ (.A1(_06217_),
    .A2(_06265_),
    .ZN(_06287_));
 NOR2_X2 _29793_ (.A1(_22508_),
    .A2(_06270_),
    .ZN(_06288_));
 AOI22_X4 _29794_ (.A1(_06271_),
    .A2(_06286_),
    .B1(_06287_),
    .B2(_06288_),
    .ZN(_06289_));
 XOR2_X1 _29795_ (.A(_06214_),
    .B(_06289_),
    .Z(_06290_));
 NOR2_X1 _29796_ (.A1(_06208_),
    .A2(_06275_),
    .ZN(_06291_));
 AOI21_X4 _29797_ (.A(_06291_),
    .B1(_06264_),
    .B2(_06209_),
    .ZN(_06292_));
 XNOR2_X2 _29798_ (.A(_06218_),
    .B(_06292_),
    .ZN(_06293_));
 XOR2_X1 _29799_ (.A(_14198_),
    .B(_22484_),
    .Z(_06294_));
 NAND2_X1 _29800_ (.A1(_06209_),
    .A2(_06294_),
    .ZN(_06295_));
 XOR2_X1 _29801_ (.A(_14202_),
    .B(_22529_),
    .Z(_06296_));
 NAND2_X1 _29802_ (.A1(_06271_),
    .A2(_06296_),
    .ZN(_06297_));
 NAND2_X4 _29803_ (.A1(_06295_),
    .A2(_06297_),
    .ZN(_06298_));
 NOR2_X2 _29804_ (.A1(_06293_),
    .A2(_06298_),
    .ZN(_06299_));
 NOR2_X2 _29805_ (.A1(_22541_),
    .A2(_06210_),
    .ZN(_06300_));
 NAND4_X4 _29806_ (.A1(_06285_),
    .A2(_06290_),
    .A3(_06299_),
    .A4(_06300_),
    .ZN(_06301_));
 INV_X1 _29807_ (.A(_00602_),
    .ZN(_06302_));
 INV_X1 _29808_ (.A(_22462_),
    .ZN(_06303_));
 MUX2_X1 _29809_ (.A(_06302_),
    .B(_06303_),
    .S(_06101_),
    .Z(_06304_));
 AOI21_X1 _29810_ (.A(_06075_),
    .B1(_06131_),
    .B2(_06304_),
    .ZN(_06305_));
 AOI211_X2 _29811_ (.A(_06126_),
    .B(_06305_),
    .C1(_06136_),
    .C2(_06127_),
    .ZN(_06306_));
 AND3_X1 _29812_ (.A1(_06177_),
    .A2(_06184_),
    .A3(_06186_),
    .ZN(_06307_));
 MUX2_X2 _29813_ (.A(_06306_),
    .B(_06307_),
    .S(_06170_),
    .Z(_06308_));
 AND4_X2 _29814_ (.A1(_06285_),
    .A2(_06290_),
    .A3(_06299_),
    .A4(_06300_),
    .ZN(_06309_));
 OAI21_X2 _29815_ (.A(_06126_),
    .B1(_06198_),
    .B2(_06199_),
    .ZN(_06310_));
 OAI21_X2 _29816_ (.A(_06309_),
    .B1(_06310_),
    .B2(_06171_),
    .ZN(_06311_));
 OAI22_X4 _29817_ (.A1(_06125_),
    .A2(_06301_),
    .B1(_06308_),
    .B2(_06311_),
    .ZN(_06312_));
 NAND3_X2 _29818_ (.A1(_06284_),
    .A2(_06290_),
    .A3(_06299_),
    .ZN(_06313_));
 OR4_X1 _29819_ (.A1(_22539_),
    .A2(_06164_),
    .A3(_06271_),
    .A4(_06313_),
    .ZN(_06314_));
 AND2_X1 _29820_ (.A1(_06074_),
    .A2(_06197_),
    .ZN(_06315_));
 MUX2_X1 _29821_ (.A(_06155_),
    .B(_06158_),
    .S(_06132_),
    .Z(_06316_));
 AOI211_X2 _29822_ (.A(_06178_),
    .B(_06315_),
    .C1(_06316_),
    .C2(_06127_),
    .ZN(_06317_));
 NAND2_X1 _29823_ (.A1(_06153_),
    .A2(_06317_),
    .ZN(_06318_));
 OAI21_X1 _29824_ (.A(_06074_),
    .B1(_06132_),
    .B2(_06137_),
    .ZN(_06319_));
 INV_X1 _29825_ (.A(_22465_),
    .ZN(_06320_));
 INV_X1 _29826_ (.A(_00603_),
    .ZN(_06321_));
 MUX2_X1 _29827_ (.A(_06320_),
    .B(_06321_),
    .S(_06101_),
    .Z(_06322_));
 INV_X1 _29828_ (.A(_00606_),
    .ZN(_06323_));
 INV_X1 _29829_ (.A(_22459_),
    .ZN(_06324_));
 MUX2_X1 _29830_ (.A(_06323_),
    .B(_06324_),
    .S(_06102_),
    .Z(_06325_));
 MUX2_X1 _29831_ (.A(_06322_),
    .B(_06325_),
    .S(_06131_),
    .Z(_06326_));
 OAI211_X2 _29832_ (.A(_06178_),
    .B(_06319_),
    .C1(_06326_),
    .C2(_06074_),
    .ZN(_06327_));
 NAND3_X1 _29833_ (.A1(_06178_),
    .A2(_06184_),
    .A3(_06186_),
    .ZN(_06328_));
 MUX2_X2 _29834_ (.A(_06327_),
    .B(_06328_),
    .S(_06171_),
    .Z(_06329_));
 AOI21_X4 _29835_ (.A(_06314_),
    .B1(_06318_),
    .B2(_06329_),
    .ZN(_06330_));
 INV_X1 _29836_ (.A(_06215_),
    .ZN(_06331_));
 OAI21_X1 _29837_ (.A(_06209_),
    .B1(_06221_),
    .B2(_06228_),
    .ZN(_06332_));
 AOI21_X1 _29838_ (.A(_06214_),
    .B1(_22501_),
    .B2(_06270_),
    .ZN(_06333_));
 NAND2_X1 _29839_ (.A1(_06332_),
    .A2(_06333_),
    .ZN(_06334_));
 OR2_X1 _29840_ (.A1(_06240_),
    .A2(_06249_),
    .ZN(_06335_));
 NOR2_X1 _29841_ (.A1(_22501_),
    .A2(_06209_),
    .ZN(_06336_));
 AOI22_X4 _29842_ (.A1(_22504_),
    .A2(_06209_),
    .B1(_06335_),
    .B2(_06336_),
    .ZN(_06337_));
 AOI21_X4 _29843_ (.A(_06331_),
    .B1(_06334_),
    .B2(_06337_),
    .ZN(_06338_));
 AND3_X2 _29844_ (.A1(_06331_),
    .A2(_06334_),
    .A3(_06337_),
    .ZN(_06339_));
 OR2_X4 _29845_ (.A1(_06338_),
    .A2(_06339_),
    .ZN(_06340_));
 XNOR2_X2 _29846_ (.A(_06214_),
    .B(_06289_),
    .ZN(_06341_));
 OR2_X1 _29847_ (.A1(_22515_),
    .A2(_22532_),
    .ZN(_06342_));
 AOI21_X1 _29848_ (.A(_06342_),
    .B1(_06226_),
    .B2(_06227_),
    .ZN(_06343_));
 AND3_X1 _29849_ (.A1(_06276_),
    .A2(_06248_),
    .A3(_06247_),
    .ZN(_06344_));
 NOR2_X1 _29850_ (.A1(_06218_),
    .A2(_06242_),
    .ZN(_06345_));
 NAND2_X1 _29851_ (.A1(_06238_),
    .A2(_06270_),
    .ZN(_06346_));
 OAI33_X1 _29852_ (.A1(_06270_),
    .A2(_06219_),
    .A3(_06343_),
    .B1(_06344_),
    .B2(_06345_),
    .B3(_06346_),
    .ZN(_06347_));
 XNOR2_X2 _29853_ (.A(_06216_),
    .B(_06347_),
    .ZN(_06348_));
 XNOR2_X2 _29854_ (.A(_06276_),
    .B(_06292_),
    .ZN(_06349_));
 NAND2_X1 _29855_ (.A1(_06209_),
    .A2(_06226_),
    .ZN(_06350_));
 OAI21_X2 _29856_ (.A(_06350_),
    .B1(_06247_),
    .B2(_06209_),
    .ZN(_06351_));
 XNOR2_X2 _29857_ (.A(_06248_),
    .B(_06351_),
    .ZN(_06352_));
 MUX2_X2 _29858_ (.A(_14203_),
    .B(_14199_),
    .S(_06210_),
    .Z(_06353_));
 NOR2_X1 _29859_ (.A1(_06298_),
    .A2(_06353_),
    .ZN(_06354_));
 OAI21_X1 _29860_ (.A(_06349_),
    .B1(_06352_),
    .B2(_06354_),
    .ZN(_06355_));
 AOI21_X2 _29861_ (.A(_06341_),
    .B1(_06348_),
    .B2(_06355_),
    .ZN(_06356_));
 OAI21_X4 _29862_ (.A(_06285_),
    .B1(_06340_),
    .B2(_06356_),
    .ZN(_06357_));
 INV_X1 _29863_ (.A(_06211_),
    .ZN(_06358_));
 OAI21_X1 _29864_ (.A(_06237_),
    .B1(_06240_),
    .B2(_06249_),
    .ZN(_06359_));
 AOI21_X1 _29865_ (.A(_06208_),
    .B1(_06280_),
    .B2(_06279_),
    .ZN(_06360_));
 AND2_X1 _29866_ (.A1(_06359_),
    .A2(_06360_),
    .ZN(_06361_));
 NOR2_X1 _29867_ (.A1(_22490_),
    .A2(_06270_),
    .ZN(_06362_));
 INV_X1 _29868_ (.A(_22487_),
    .ZN(_06363_));
 NOR2_X1 _29869_ (.A1(_06363_),
    .A2(_06208_),
    .ZN(_06364_));
 OR2_X1 _29870_ (.A1(_06362_),
    .A2(_06364_),
    .ZN(_06365_));
 NAND2_X1 _29871_ (.A1(_06213_),
    .A2(_06211_),
    .ZN(_06366_));
 NOR3_X1 _29872_ (.A1(_06270_),
    .A2(_06229_),
    .A3(_06232_),
    .ZN(_06367_));
 OAI33_X1 _29873_ (.A1(_06358_),
    .A2(_06361_),
    .A3(_06365_),
    .B1(_06366_),
    .B2(_06367_),
    .B3(_06364_),
    .ZN(_06368_));
 AOI21_X1 _29874_ (.A(_06365_),
    .B1(_06360_),
    .B2(_06359_),
    .ZN(_06369_));
 NOR2_X1 _29875_ (.A1(_06212_),
    .A2(_06364_),
    .ZN(_06370_));
 OR3_X1 _29876_ (.A1(_06270_),
    .A2(_06229_),
    .A3(_06232_),
    .ZN(_06371_));
 AOI211_X2 _29877_ (.A(_06211_),
    .B(_06369_),
    .C1(_06370_),
    .C2(_06371_),
    .ZN(_06372_));
 NOR2_X4 _29878_ (.A1(net342),
    .A2(_06372_),
    .ZN(_06373_));
 NAND2_X2 _29879_ (.A1(_06357_),
    .A2(_06373_),
    .ZN(_06374_));
 NOR4_X4 _29880_ (.A1(_06258_),
    .A2(_06312_),
    .A3(_06330_),
    .A4(_06374_),
    .ZN(_06375_));
 BUF_X4 _29881_ (.A(_06258_),
    .Z(_06376_));
 NOR3_X4 _29882_ (.A1(_06165_),
    .A2(_06171_),
    .A3(_06256_),
    .ZN(_06377_));
 NAND2_X1 _29883_ (.A1(_22497_),
    .A2(_06210_),
    .ZN(_06378_));
 NAND3_X2 _29884_ (.A1(_06254_),
    .A2(_06363_),
    .A3(_06271_),
    .ZN(_06379_));
 AND3_X1 _29885_ (.A1(_06212_),
    .A2(_06281_),
    .A3(_06278_),
    .ZN(_06380_));
 OAI21_X4 _29886_ (.A(_06378_),
    .B1(_06379_),
    .B2(_06380_),
    .ZN(_06381_));
 NAND3_X1 _29887_ (.A1(_06213_),
    .A2(_06260_),
    .A3(_06266_),
    .ZN(_06382_));
 AOI221_X2 _29888_ (.A(_06211_),
    .B1(_22494_),
    .B2(_06271_),
    .C1(_06382_),
    .C2(_06362_),
    .ZN(_06383_));
 NOR2_X4 _29889_ (.A1(_06381_),
    .A2(_06383_),
    .ZN(_06384_));
 XNOR2_X2 _29890_ (.A(_06377_),
    .B(_06384_),
    .ZN(_06385_));
 CLKBUF_X3 _29891_ (.A(_06385_),
    .Z(_06386_));
 NOR2_X2 _29892_ (.A1(_06376_),
    .A2(_06386_),
    .ZN(_06387_));
 OR2_X1 _29893_ (.A1(_06375_),
    .A2(_06387_),
    .ZN(_22545_));
 BUF_X2 _29894_ (.A(_22548_),
    .Z(_06388_));
 NOR4_X4 _29895_ (.A1(_06338_),
    .A2(_06339_),
    .A3(_06368_),
    .A4(_06372_),
    .ZN(_06389_));
 OR4_X4 _29896_ (.A1(_06267_),
    .A2(_06269_),
    .A3(_06282_),
    .A4(_06283_),
    .ZN(_06390_));
 AND2_X1 _29897_ (.A1(_06295_),
    .A2(_06297_),
    .ZN(_06391_));
 XNOR2_X2 _29898_ (.A(_06227_),
    .B(_06351_),
    .ZN(_06392_));
 AND4_X2 _29899_ (.A1(_06349_),
    .A2(_06391_),
    .A3(_06348_),
    .A4(_06392_),
    .ZN(_06393_));
 NOR3_X2 _29900_ (.A1(_06390_),
    .A2(_06341_),
    .A3(_06393_),
    .ZN(_06394_));
 OR2_X1 _29901_ (.A1(_06253_),
    .A2(_06381_),
    .ZN(_06395_));
 AOI221_X1 _29902_ (.A(_06210_),
    .B1(_06389_),
    .B2(_06394_),
    .C1(_06395_),
    .C2(_06254_),
    .ZN(_06396_));
 OR2_X1 _29903_ (.A1(_22497_),
    .A2(_06235_),
    .ZN(_06397_));
 AOI221_X1 _29904_ (.A(_06384_),
    .B1(_06389_),
    .B2(_06394_),
    .C1(_06397_),
    .C2(_06210_),
    .ZN(_06398_));
 OR3_X1 _29905_ (.A1(_06165_),
    .A2(_06171_),
    .A3(_06256_),
    .ZN(_06399_));
 BUF_X4 _29906_ (.A(_06399_),
    .Z(_06400_));
 MUX2_X1 _29907_ (.A(_06396_),
    .B(_06398_),
    .S(_06400_),
    .Z(_06401_));
 XNOR2_X2 _29908_ (.A(_06388_),
    .B(_06401_),
    .ZN(_06402_));
 INV_X2 _29909_ (.A(_06402_),
    .ZN(_19434_));
 BUF_X1 _29910_ (.A(_14209_),
    .Z(_06403_));
 INV_X1 _29911_ (.A(_06403_),
    .ZN(_06404_));
 BUF_X4 _29912_ (.A(_06404_),
    .Z(_06405_));
 BUF_X4 _29913_ (.A(_06405_),
    .Z(_14204_));
 XNOR2_X2 _29914_ (.A(_06400_),
    .B(_06384_),
    .ZN(_06406_));
 BUF_X4 _29915_ (.A(_06406_),
    .Z(_06407_));
 NOR2_X4 _29916_ (.A1(_06338_),
    .A2(_06339_),
    .ZN(_06408_));
 INV_X1 _29917_ (.A(_06348_),
    .ZN(_06409_));
 AND2_X1 _29918_ (.A1(_14199_),
    .A2(_06210_),
    .ZN(_06410_));
 AOI21_X4 _29919_ (.A(_06410_),
    .B1(_06271_),
    .B2(_14203_),
    .ZN(_06411_));
 NAND2_X1 _29920_ (.A1(_06391_),
    .A2(_06411_),
    .ZN(_06412_));
 AOI21_X1 _29921_ (.A(_06293_),
    .B1(_06392_),
    .B2(_06412_),
    .ZN(_06413_));
 OAI21_X2 _29922_ (.A(_06290_),
    .B1(_06409_),
    .B2(_06413_),
    .ZN(_06414_));
 AOI21_X4 _29923_ (.A(_06390_),
    .B1(_06408_),
    .B2(_06414_),
    .ZN(_06415_));
 OR2_X1 _29924_ (.A1(_06368_),
    .A2(_06372_),
    .ZN(_06416_));
 CLKBUF_X3 _29925_ (.A(_06416_),
    .Z(_06417_));
 NOR2_X4 _29926_ (.A1(_06415_),
    .A2(_06417_),
    .ZN(_06418_));
 NOR4_X2 _29927_ (.A1(_14204_),
    .A2(_06376_),
    .A3(_06407_),
    .A4(_06418_),
    .ZN(_06419_));
 CLKBUF_X3 _29928_ (.A(_22544_),
    .Z(_06420_));
 INV_X1 _29929_ (.A(_06420_),
    .ZN(_06421_));
 BUF_X4 _29930_ (.A(_06271_),
    .Z(_06422_));
 AOI21_X1 _29931_ (.A(_06422_),
    .B1(_06317_),
    .B2(_06153_),
    .ZN(_06423_));
 NOR2_X1 _29932_ (.A1(_06165_),
    .A2(_06210_),
    .ZN(_06424_));
 MUX2_X2 _29933_ (.A(_06423_),
    .B(_06424_),
    .S(_06308_),
    .Z(_06425_));
 NAND4_X2 _29934_ (.A1(_06125_),
    .A2(_06153_),
    .A3(_06422_),
    .A4(_06317_),
    .ZN(_06426_));
 OAI21_X4 _29935_ (.A(_06426_),
    .B1(_06422_),
    .B2(_06125_),
    .ZN(_06427_));
 OAI21_X1 _29936_ (.A(_06421_),
    .B1(_06425_),
    .B2(_06427_),
    .ZN(_06428_));
 OAI21_X1 _29937_ (.A(_06254_),
    .B1(_06253_),
    .B2(_06381_),
    .ZN(_06429_));
 NAND2_X1 _29938_ (.A1(_06422_),
    .A2(_06429_),
    .ZN(_06430_));
 OR2_X2 _29939_ (.A1(_06381_),
    .A2(_06383_),
    .ZN(_06431_));
 NAND2_X1 _29940_ (.A1(_06236_),
    .A2(_06431_),
    .ZN(_06432_));
 MUX2_X2 _29941_ (.A(_06430_),
    .B(_06432_),
    .S(_06400_),
    .Z(_06433_));
 INV_X1 _29942_ (.A(_22539_),
    .ZN(_06434_));
 INV_X1 _29943_ (.A(_22541_),
    .ZN(_06435_));
 MUX2_X2 _29944_ (.A(_06434_),
    .B(_06435_),
    .S(_06422_),
    .Z(_06436_));
 OAI21_X1 _29945_ (.A(_06433_),
    .B1(_06436_),
    .B2(_06353_),
    .ZN(_06437_));
 OAI22_X2 _29946_ (.A1(_06419_),
    .A2(_06428_),
    .B1(_06437_),
    .B2(_06421_),
    .ZN(_06438_));
 NAND3_X1 _29947_ (.A1(_06403_),
    .A2(_06407_),
    .A3(_06436_),
    .ZN(_06439_));
 NOR3_X1 _29948_ (.A1(_06405_),
    .A2(_06165_),
    .A3(_06422_),
    .ZN(_06440_));
 NOR2_X2 _29949_ (.A1(_06171_),
    .A2(_06310_),
    .ZN(_06441_));
 OAI21_X1 _29950_ (.A(_06440_),
    .B1(_06441_),
    .B2(_06308_),
    .ZN(_06442_));
 NAND2_X1 _29951_ (.A1(_06403_),
    .A2(_06422_),
    .ZN(_06443_));
 OR3_X1 _29952_ (.A1(_06308_),
    .A2(_06441_),
    .A3(_06443_),
    .ZN(_06444_));
 OR2_X1 _29953_ (.A1(_06125_),
    .A2(_06443_),
    .ZN(_06445_));
 NAND4_X1 _29954_ (.A1(_06386_),
    .A2(_06442_),
    .A3(_06444_),
    .A4(_06445_),
    .ZN(_06446_));
 NOR3_X2 _29955_ (.A1(_06312_),
    .A2(_06330_),
    .A3(_06374_),
    .ZN(_06447_));
 AOI21_X2 _29956_ (.A(_06301_),
    .B1(_06317_),
    .B2(_06153_),
    .ZN(_06448_));
 AOI22_X4 _29957_ (.A1(_06165_),
    .A2(_06309_),
    .B1(_06329_),
    .B2(_06448_),
    .ZN(_06449_));
 NOR4_X4 _29958_ (.A1(_22539_),
    .A2(_06165_),
    .A3(_06422_),
    .A4(_06313_),
    .ZN(_06450_));
 OAI21_X4 _29959_ (.A(_06450_),
    .B1(_06441_),
    .B2(_06308_),
    .ZN(_06451_));
 NAND2_X1 _29960_ (.A1(_06449_),
    .A2(_06451_),
    .ZN(_06452_));
 CLKBUF_X3 _29961_ (.A(_06373_),
    .Z(_06453_));
 NAND4_X2 _29962_ (.A1(_06403_),
    .A2(_06357_),
    .A3(_06453_),
    .A4(_06436_),
    .ZN(_06454_));
 OAI221_X2 _29963_ (.A(_06439_),
    .B1(_06446_),
    .B2(_06447_),
    .C1(_06452_),
    .C2(_06454_),
    .ZN(_06455_));
 CLKBUF_X3 _29964_ (.A(_06433_),
    .Z(_06456_));
 MUX2_X2 _29965_ (.A(_22539_),
    .B(_22541_),
    .S(_06422_),
    .Z(_06457_));
 OAI21_X1 _29966_ (.A(_06456_),
    .B1(_06457_),
    .B2(_06420_),
    .ZN(_06458_));
 NOR2_X1 _29967_ (.A1(_06405_),
    .A2(_06376_),
    .ZN(_06459_));
 OAI22_X4 _29968_ (.A1(_06407_),
    .A2(_06418_),
    .B1(_06425_),
    .B2(_06427_),
    .ZN(_06460_));
 NAND2_X1 _29969_ (.A1(_06459_),
    .A2(_06460_),
    .ZN(_06461_));
 AND2_X1 _29970_ (.A1(_06400_),
    .A2(_06432_),
    .ZN(_06462_));
 AOI21_X4 _29971_ (.A(_06462_),
    .B1(_06430_),
    .B2(_06377_),
    .ZN(_06463_));
 BUF_X4 _29972_ (.A(_06463_),
    .Z(_06464_));
 AOI221_X2 _29973_ (.A(_06438_),
    .B1(_06455_),
    .B2(_06458_),
    .C1(_06461_),
    .C2(_06464_),
    .ZN(_06465_));
 INV_X1 _29974_ (.A(_06465_),
    .ZN(_06466_));
 NOR2_X2 _29975_ (.A1(_06390_),
    .A2(_06341_),
    .ZN(_06467_));
 AND2_X2 _29976_ (.A1(_06467_),
    .A2(_06389_),
    .ZN(_06468_));
 NAND3_X1 _29977_ (.A1(_14199_),
    .A2(_06434_),
    .A3(_06210_),
    .ZN(_06469_));
 NAND3_X1 _29978_ (.A1(_14203_),
    .A2(_06435_),
    .A3(_06271_),
    .ZN(_06470_));
 NAND3_X1 _29979_ (.A1(_06391_),
    .A2(_06469_),
    .A3(_06470_),
    .ZN(_06471_));
 OAI21_X1 _29980_ (.A(_06349_),
    .B1(_06352_),
    .B2(_06471_),
    .ZN(_06472_));
 OAI21_X2 _29981_ (.A(_06290_),
    .B1(_06409_),
    .B2(_06472_),
    .ZN(_06473_));
 OAI211_X4 _29982_ (.A(_06285_),
    .B(_06373_),
    .C1(_06473_),
    .C2(_06340_),
    .ZN(_06474_));
 NOR2_X1 _29983_ (.A1(_06415_),
    .A2(_06474_),
    .ZN(_06475_));
 NAND4_X4 _29984_ (.A1(_06449_),
    .A2(_06451_),
    .A3(_06468_),
    .A4(_06475_),
    .ZN(_06476_));
 AOI21_X4 _29985_ (.A(_06433_),
    .B1(_06468_),
    .B2(_06393_),
    .ZN(_06477_));
 NAND3_X2 _29986_ (.A1(_19434_),
    .A2(_06476_),
    .A3(_06477_),
    .ZN(_06478_));
 NOR3_X1 _29987_ (.A1(_06425_),
    .A2(_06427_),
    .A3(_06436_),
    .ZN(_06479_));
 OAI21_X1 _29988_ (.A(_06456_),
    .B1(_06479_),
    .B2(_06420_),
    .ZN(_06480_));
 AOI21_X1 _29989_ (.A(_06466_),
    .B1(_06478_),
    .B2(_06480_),
    .ZN(_22551_));
 CLKBUF_X3 _29990_ (.A(_06061_),
    .Z(_06481_));
 NOR2_X1 _29991_ (.A1(\g_reduce0[14].adder.x[0] ),
    .A2(_06481_),
    .ZN(_06482_));
 NOR4_X4 _29992_ (.A1(_06057_),
    .A2(_06058_),
    .A3(_06059_),
    .A4(_06060_),
    .ZN(_06483_));
 AOI21_X1 _29993_ (.A(_06483_),
    .B1(_06064_),
    .B2(\g_reduce0[12].adder.x[0] ),
    .ZN(_06484_));
 OR4_X4 _29994_ (.A1(\g_reduce0[14].adder.x[11] ),
    .A2(\g_reduce0[14].adder.x[12] ),
    .A3(_06062_),
    .A4(_06063_),
    .ZN(_06485_));
 BUF_X4 _29995_ (.A(_06485_),
    .Z(_06486_));
 NAND2_X1 _29996_ (.A1(_06456_),
    .A2(_06428_),
    .ZN(_06487_));
 OAI21_X1 _29997_ (.A(_06487_),
    .B1(_06478_),
    .B2(_06461_),
    .ZN(_06488_));
 NAND2_X1 _29998_ (.A1(_06420_),
    .A2(_06456_),
    .ZN(_06489_));
 OAI21_X1 _29999_ (.A(_06488_),
    .B1(_06489_),
    .B2(_06457_),
    .ZN(_06490_));
 OR2_X1 _30000_ (.A1(_06415_),
    .A2(_06474_),
    .ZN(_06491_));
 NAND4_X1 _30001_ (.A1(_06422_),
    .A2(_06467_),
    .A3(_06389_),
    .A4(_06429_),
    .ZN(_06492_));
 NAND4_X1 _30002_ (.A1(_06236_),
    .A2(_06431_),
    .A3(_06467_),
    .A4(_06389_),
    .ZN(_06493_));
 MUX2_X2 _30003_ (.A(_06492_),
    .B(_06493_),
    .S(_06400_),
    .Z(_06494_));
 NOR4_X4 _30004_ (.A1(_06312_),
    .A2(_06330_),
    .A3(_06491_),
    .A4(_06494_),
    .ZN(_06495_));
 AND2_X2 _30005_ (.A1(_06389_),
    .A2(_06394_),
    .ZN(_06496_));
 NOR2_X2 _30006_ (.A1(_06496_),
    .A2(_06494_),
    .ZN(_06497_));
 NOR3_X4 _30007_ (.A1(_06376_),
    .A2(_06495_),
    .A3(_06497_),
    .ZN(_19438_));
 NAND3_X1 _30008_ (.A1(_22546_),
    .A2(_19434_),
    .A3(_19438_),
    .ZN(_06498_));
 BUF_X4 _30009_ (.A(_06464_),
    .Z(_06499_));
 AOI21_X1 _30010_ (.A(_06490_),
    .B1(_06498_),
    .B2(_06499_),
    .ZN(_06500_));
 OAI21_X1 _30011_ (.A(_06458_),
    .B1(_06478_),
    .B2(_06455_),
    .ZN(_06501_));
 OAI21_X1 _30012_ (.A(_06501_),
    .B1(_06489_),
    .B2(_06411_),
    .ZN(_06502_));
 MUX2_X1 _30013_ (.A(_06490_),
    .B(_06500_),
    .S(_06502_),
    .Z(_06503_));
 AND2_X1 _30014_ (.A1(_06476_),
    .A2(_06477_),
    .ZN(_06504_));
 CLKBUF_X3 _30015_ (.A(_06402_),
    .Z(_06505_));
 AND2_X1 _30016_ (.A1(_06236_),
    .A2(_06257_),
    .ZN(_06506_));
 CLKBUF_X3 _30017_ (.A(_06506_),
    .Z(_06507_));
 NAND2_X1 _30018_ (.A1(_06403_),
    .A2(_06507_),
    .ZN(_06508_));
 NAND2_X1 _30019_ (.A1(_06386_),
    .A2(_06417_),
    .ZN(_06509_));
 AOI21_X1 _30020_ (.A(_06341_),
    .B1(_06453_),
    .B2(_06390_),
    .ZN(_06510_));
 AOI221_X2 _30021_ (.A(_06508_),
    .B1(_06509_),
    .B2(_06408_),
    .C1(_06510_),
    .C2(_06386_),
    .ZN(_06511_));
 NAND2_X1 _30022_ (.A1(_06505_),
    .A2(_06511_),
    .ZN(_06512_));
 NOR3_X1 _30023_ (.A1(_06285_),
    .A2(_06453_),
    .A3(_06505_),
    .ZN(_06513_));
 NOR2_X1 _30024_ (.A1(_06341_),
    .A2(_06348_),
    .ZN(_06514_));
 OAI21_X1 _30025_ (.A(_06285_),
    .B1(_06340_),
    .B2(_06514_),
    .ZN(_06515_));
 NAND2_X1 _30026_ (.A1(_06373_),
    .A2(_06515_),
    .ZN(_06516_));
 AOI211_X2 _30027_ (.A(_06258_),
    .B(_06348_),
    .C1(_06516_),
    .C2(_06386_),
    .ZN(_06517_));
 NOR2_X1 _30028_ (.A1(_06384_),
    .A2(_06373_),
    .ZN(_06518_));
 NOR2_X1 _30029_ (.A1(_06431_),
    .A2(_06373_),
    .ZN(_06519_));
 MUX2_X1 _30030_ (.A(_06518_),
    .B(_06519_),
    .S(_06377_),
    .Z(_06520_));
 AND3_X1 _30031_ (.A1(_06507_),
    .A2(_06293_),
    .A3(_06520_),
    .ZN(_06521_));
 NOR3_X1 _30032_ (.A1(_06349_),
    .A2(_06433_),
    .A3(_06515_),
    .ZN(_06522_));
 OR3_X1 _30033_ (.A1(_06517_),
    .A2(_06521_),
    .A3(_06522_),
    .ZN(_06523_));
 AOI21_X1 _30034_ (.A(_06513_),
    .B1(_06523_),
    .B2(_06505_),
    .ZN(_06524_));
 CLKBUF_X3 _30035_ (.A(_06403_),
    .Z(_06525_));
 OAI21_X1 _30036_ (.A(_06512_),
    .B1(_06524_),
    .B2(_06525_),
    .ZN(_06526_));
 AND2_X1 _30037_ (.A1(_06504_),
    .A2(_06526_),
    .ZN(_06527_));
 AND2_X1 _30038_ (.A1(_06459_),
    .A2(_06460_),
    .ZN(_06528_));
 NAND2_X1 _30039_ (.A1(_06505_),
    .A2(_06528_),
    .ZN(_06529_));
 NOR4_X2 _30040_ (.A1(_06376_),
    .A2(_06353_),
    .A3(_06415_),
    .A4(_06417_),
    .ZN(_06530_));
 NOR2_X1 _30041_ (.A1(_06373_),
    .A2(_06436_),
    .ZN(_06531_));
 MUX2_X1 _30042_ (.A(_06411_),
    .B(_06531_),
    .S(_06385_),
    .Z(_06532_));
 NAND3_X2 _30043_ (.A1(_06449_),
    .A2(_06451_),
    .A3(_06357_),
    .ZN(_06533_));
 NOR2_X1 _30044_ (.A1(_06433_),
    .A2(_06436_),
    .ZN(_06534_));
 AOI221_X2 _30045_ (.A(_06530_),
    .B1(_06532_),
    .B2(_06507_),
    .C1(_06533_),
    .C2(_06534_),
    .ZN(_06535_));
 NAND3_X1 _30046_ (.A1(_06236_),
    .A2(_06257_),
    .A3(_06298_),
    .ZN(_06536_));
 OAI33_X1 _30047_ (.A1(_06391_),
    .A2(_06357_),
    .A3(_06433_),
    .B1(_06536_),
    .B2(_06453_),
    .B3(_06407_),
    .ZN(_06537_));
 BUF_X2 _30048_ (.A(_06386_),
    .Z(_06538_));
 NAND2_X1 _30049_ (.A1(_06293_),
    .A2(_06348_),
    .ZN(_06539_));
 AOI21_X1 _30050_ (.A(_06340_),
    .B1(_06539_),
    .B2(_06290_),
    .ZN(_06540_));
 OAI21_X1 _30051_ (.A(_06453_),
    .B1(_06540_),
    .B2(_06390_),
    .ZN(_06541_));
 AOI21_X1 _30052_ (.A(_06376_),
    .B1(_06538_),
    .B2(_06541_),
    .ZN(_06542_));
 AOI21_X2 _30053_ (.A(_06537_),
    .B1(_06542_),
    .B2(_06352_),
    .ZN(_06543_));
 MUX2_X2 _30054_ (.A(_06535_),
    .B(_06543_),
    .S(_06525_),
    .Z(_06544_));
 OAI21_X1 _30055_ (.A(_06529_),
    .B1(_06544_),
    .B2(_06505_),
    .ZN(_06545_));
 OR2_X1 _30056_ (.A1(_06495_),
    .A2(_06497_),
    .ZN(_06546_));
 CLKBUF_X3 _30057_ (.A(_06421_),
    .Z(_06547_));
 AOI221_X2 _30058_ (.A(_06527_),
    .B1(_06545_),
    .B2(_06546_),
    .C1(_06376_),
    .C2(_06547_),
    .ZN(_06548_));
 BUF_X2 _30059_ (.A(_06548_),
    .Z(_06549_));
 MUX2_X1 _30060_ (.A(_06285_),
    .B(_06453_),
    .S(_06420_),
    .Z(_06550_));
 NOR2_X1 _30061_ (.A1(_06464_),
    .A2(_06550_),
    .ZN(_06551_));
 OAI221_X2 _30062_ (.A(_06405_),
    .B1(_06506_),
    .B2(_06353_),
    .C1(_06536_),
    .C2(_06385_),
    .ZN(_06552_));
 NOR2_X1 _30063_ (.A1(_06407_),
    .A2(_06353_),
    .ZN(_06553_));
 NAND3_X2 _30064_ (.A1(_06449_),
    .A2(_06451_),
    .A3(_06418_),
    .ZN(_06554_));
 AOI221_X2 _30065_ (.A(_06552_),
    .B1(_06553_),
    .B2(_06554_),
    .C1(_06298_),
    .C2(_06375_),
    .ZN(_06555_));
 NAND3_X2 _30066_ (.A1(_06505_),
    .A2(_06476_),
    .A3(_06477_),
    .ZN(_06556_));
 NAND4_X1 _30067_ (.A1(_06506_),
    .A2(_06449_),
    .A3(_06451_),
    .A4(_06418_),
    .ZN(_06557_));
 AOI21_X1 _30068_ (.A(_06392_),
    .B1(_06406_),
    .B2(_06506_),
    .ZN(_06558_));
 AOI21_X1 _30069_ (.A(_06258_),
    .B1(_06386_),
    .B2(_06516_),
    .ZN(_06559_));
 AOI221_X2 _30070_ (.A(_06405_),
    .B1(_06557_),
    .B2(_06558_),
    .C1(_06559_),
    .C2(_06293_),
    .ZN(_06560_));
 NOR3_X1 _30071_ (.A1(_06555_),
    .A2(_06556_),
    .A3(_06560_),
    .ZN(_06561_));
 NOR2_X1 _30072_ (.A1(_06525_),
    .A2(_06290_),
    .ZN(_06562_));
 OAI21_X1 _30073_ (.A(_06562_),
    .B1(_06447_),
    .B2(_06407_),
    .ZN(_06563_));
 NOR2_X1 _30074_ (.A1(_06400_),
    .A2(_06384_),
    .ZN(_06564_));
 NOR2_X1 _30075_ (.A1(_06377_),
    .A2(_06431_),
    .ZN(_06565_));
 AND2_X1 _30076_ (.A1(_06400_),
    .A2(_06518_),
    .ZN(_06566_));
 AND2_X1 _30077_ (.A1(_06377_),
    .A2(_06519_),
    .ZN(_06567_));
 OAI33_X1 _30078_ (.A1(_06564_),
    .A2(_06565_),
    .A3(_06408_),
    .B1(_06566_),
    .B2(_06567_),
    .B3(_06285_),
    .ZN(_06568_));
 NOR3_X1 _30079_ (.A1(_06525_),
    .A2(_06407_),
    .A3(_06348_),
    .ZN(_06569_));
 AOI22_X1 _30080_ (.A1(_06525_),
    .A2(_06568_),
    .B1(_06569_),
    .B2(_06554_),
    .ZN(_06570_));
 AOI21_X1 _30081_ (.A(_06478_),
    .B1(_06563_),
    .B2(_06570_),
    .ZN(_06571_));
 NAND2_X1 _30082_ (.A1(_06389_),
    .A2(_06394_),
    .ZN(_06572_));
 NOR2_X1 _30083_ (.A1(_06572_),
    .A2(_06474_),
    .ZN(_06573_));
 OAI221_X2 _30084_ (.A(_06388_),
    .B1(_06375_),
    .B2(_06387_),
    .C1(_06456_),
    .C2(_06573_),
    .ZN(_06574_));
 OR2_X1 _30085_ (.A1(_06388_),
    .A2(_06496_),
    .ZN(_06575_));
 AOI211_X2 _30086_ (.A(_06455_),
    .B(_06494_),
    .C1(_06574_),
    .C2(_06575_),
    .ZN(_06576_));
 OR4_X2 _30087_ (.A1(_06551_),
    .A2(_06561_),
    .A3(_06571_),
    .A4(_06576_),
    .ZN(_06577_));
 XNOR2_X2 _30088_ (.A(_06388_),
    .B(_06496_),
    .ZN(_06578_));
 NAND2_X2 _30089_ (.A1(_06463_),
    .A2(_06578_),
    .ZN(_06579_));
 AOI221_X2 _30090_ (.A(_06511_),
    .B1(_06546_),
    .B2(_06528_),
    .C1(_06523_),
    .C2(_14204_),
    .ZN(_06580_));
 MUX2_X1 _30091_ (.A(_06285_),
    .B(_06408_),
    .S(_06547_),
    .Z(_06581_));
 OAI222_X2 _30092_ (.A1(_06544_),
    .A2(_06556_),
    .B1(_06579_),
    .B2(_06580_),
    .C1(_06581_),
    .C2(_06464_),
    .ZN(_06582_));
 MUX2_X1 _30093_ (.A(_06341_),
    .B(_06340_),
    .S(_06420_),
    .Z(_06583_));
 INV_X1 _30094_ (.A(_22546_),
    .ZN(_06584_));
 OAI21_X1 _30095_ (.A(_06463_),
    .B1(_06505_),
    .B2(_06584_),
    .ZN(_06585_));
 OAI22_X1 _30096_ (.A1(_06464_),
    .A2(_06583_),
    .B1(_06585_),
    .B2(_19438_),
    .ZN(_06586_));
 NAND3_X1 _30097_ (.A1(_14204_),
    .A2(_06507_),
    .A3(_06457_),
    .ZN(_06587_));
 AOI21_X2 _30098_ (.A(_06587_),
    .B1(_06554_),
    .B2(_06538_),
    .ZN(_06588_));
 NOR4_X1 _30099_ (.A1(_06403_),
    .A2(_06376_),
    .A3(_06425_),
    .A4(_06427_),
    .ZN(_06589_));
 AND3_X1 _30100_ (.A1(_06538_),
    .A2(_06554_),
    .A3(_06589_),
    .ZN(_06590_));
 NOR3_X1 _30101_ (.A1(_06391_),
    .A2(_06415_),
    .A3(_06417_),
    .ZN(_06591_));
 NAND3_X1 _30102_ (.A1(_06525_),
    .A2(_06507_),
    .A3(_06591_),
    .ZN(_06592_));
 AOI22_X2 _30103_ (.A1(_06407_),
    .A2(_06298_),
    .B1(_06411_),
    .B2(_06520_),
    .ZN(_06593_));
 NAND4_X1 _30104_ (.A1(_06525_),
    .A2(_06507_),
    .A3(_06386_),
    .A4(_06411_),
    .ZN(_06594_));
 NOR3_X1 _30105_ (.A1(_06312_),
    .A2(_06330_),
    .A3(_06415_),
    .ZN(_06595_));
 OAI221_X2 _30106_ (.A(_06592_),
    .B1(_06593_),
    .B2(_06508_),
    .C1(_06594_),
    .C2(_06595_),
    .ZN(_06596_));
 NOR3_X1 _30107_ (.A1(_06588_),
    .A2(_06590_),
    .A3(_06596_),
    .ZN(_06597_));
 AND3_X1 _30108_ (.A1(_06402_),
    .A2(_06476_),
    .A3(_06477_),
    .ZN(_06598_));
 NAND2_X1 _30109_ (.A1(_06476_),
    .A2(_06477_),
    .ZN(_06599_));
 NOR2_X1 _30110_ (.A1(_06505_),
    .A2(_06599_),
    .ZN(_06600_));
 OR4_X1 _30111_ (.A1(_14204_),
    .A2(_06409_),
    .A3(_06375_),
    .A4(_06387_),
    .ZN(_06601_));
 NOR2_X1 _30112_ (.A1(_14204_),
    .A2(_06341_),
    .ZN(_06602_));
 OAI21_X1 _30113_ (.A(_06602_),
    .B1(_06387_),
    .B2(_06375_),
    .ZN(_06603_));
 AND2_X1 _30114_ (.A1(_06538_),
    .A2(_06516_),
    .ZN(_06604_));
 NAND2_X1 _30115_ (.A1(_06507_),
    .A2(_06293_),
    .ZN(_06605_));
 OAI21_X1 _30116_ (.A(_06352_),
    .B1(_06538_),
    .B2(_06376_),
    .ZN(_06606_));
 OAI221_X2 _30117_ (.A(_14204_),
    .B1(_06604_),
    .B2(_06605_),
    .C1(_06606_),
    .C2(_06375_),
    .ZN(_06607_));
 NAND4_X1 _30118_ (.A1(_06507_),
    .A2(_06601_),
    .A3(_06603_),
    .A4(_06607_),
    .ZN(_06608_));
 AOI221_X4 _30119_ (.A(_06586_),
    .B1(_06597_),
    .B2(_06598_),
    .C1(_06600_),
    .C2(_06608_),
    .ZN(_06609_));
 NOR3_X1 _30120_ (.A1(_06517_),
    .A2(_06521_),
    .A3(_06522_),
    .ZN(_06610_));
 MUX2_X1 _30121_ (.A(_06610_),
    .B(_06543_),
    .S(_14204_),
    .Z(_06611_));
 NOR3_X1 _30122_ (.A1(_06405_),
    .A2(_06353_),
    .A3(_06417_),
    .ZN(_06612_));
 NAND3_X1 _30123_ (.A1(_06236_),
    .A2(_06257_),
    .A3(_06612_),
    .ZN(_06613_));
 NOR4_X2 _30124_ (.A1(_06312_),
    .A2(_06330_),
    .A3(_06415_),
    .A4(_06613_),
    .ZN(_06614_));
 OAI221_X2 _30125_ (.A(_06405_),
    .B1(_06407_),
    .B2(_06418_),
    .C1(_06425_),
    .C2(_06427_),
    .ZN(_06615_));
 OAI21_X1 _30126_ (.A(_06403_),
    .B1(_06381_),
    .B2(_06383_),
    .ZN(_06616_));
 AOI21_X1 _30127_ (.A(_06616_),
    .B1(_06457_),
    .B2(_06417_),
    .ZN(_06617_));
 OR3_X1 _30128_ (.A1(_06404_),
    .A2(_06381_),
    .A3(_06383_),
    .ZN(_06618_));
 AOI21_X1 _30129_ (.A(_06618_),
    .B1(_06457_),
    .B2(_06417_),
    .ZN(_06619_));
 MUX2_X1 _30130_ (.A(_06617_),
    .B(_06619_),
    .S(_06377_),
    .Z(_06620_));
 NOR4_X2 _30131_ (.A1(_06405_),
    .A2(_06400_),
    .A3(_06384_),
    .A4(_06411_),
    .ZN(_06621_));
 NOR4_X2 _30132_ (.A1(_06405_),
    .A2(_06377_),
    .A3(_06431_),
    .A4(_06411_),
    .ZN(_06622_));
 NOR4_X2 _30133_ (.A1(_06376_),
    .A2(_06620_),
    .A3(_06621_),
    .A4(_06622_),
    .ZN(_06623_));
 NOR3_X1 _30134_ (.A1(_06405_),
    .A2(_06433_),
    .A3(_06436_),
    .ZN(_06624_));
 AOI221_X2 _30135_ (.A(_06614_),
    .B1(_06615_),
    .B2(_06623_),
    .C1(_06624_),
    .C2(_06533_),
    .ZN(_06625_));
 AOI21_X1 _30136_ (.A(_06453_),
    .B1(_06285_),
    .B2(_06538_),
    .ZN(_06626_));
 NAND2_X1 _30137_ (.A1(_06290_),
    .A2(_06417_),
    .ZN(_06627_));
 MUX2_X1 _30138_ (.A(_06340_),
    .B(_06627_),
    .S(_06538_),
    .Z(_06628_));
 AOI221_X1 _30139_ (.A(_06403_),
    .B1(_06386_),
    .B2(_06467_),
    .C1(_06408_),
    .C2(_06453_),
    .ZN(_06629_));
 AOI22_X1 _30140_ (.A1(_06525_),
    .A2(_06626_),
    .B1(_06628_),
    .B2(_06629_),
    .ZN(_06630_));
 MUX2_X1 _30141_ (.A(_06625_),
    .B(_06630_),
    .S(_19438_),
    .Z(_06631_));
 MUX2_X1 _30142_ (.A(_06538_),
    .B(_06453_),
    .S(_06547_),
    .Z(_06632_));
 OAI222_X2 _30143_ (.A1(_06556_),
    .A2(_06611_),
    .B1(_06631_),
    .B2(_06579_),
    .C1(_06632_),
    .C2(_06499_),
    .ZN(_06633_));
 NAND4_X2 _30144_ (.A1(_06577_),
    .A2(_06582_),
    .A3(_06609_),
    .A4(_06633_),
    .ZN(_06634_));
 NAND3_X1 _30145_ (.A1(_06601_),
    .A2(_06603_),
    .A3(_06607_),
    .ZN(_06635_));
 OR2_X1 _30146_ (.A1(_06556_),
    .A2(_06635_),
    .ZN(_06636_));
 NOR2_X1 _30147_ (.A1(_06547_),
    .A2(_06507_),
    .ZN(_06637_));
 NAND2_X1 _30148_ (.A1(_06538_),
    .A2(_06453_),
    .ZN(_06638_));
 MUX2_X1 _30149_ (.A(_06568_),
    .B(_06638_),
    .S(_06525_),
    .Z(_06639_));
 AOI221_X1 _30150_ (.A(_06637_),
    .B1(_06639_),
    .B2(_06600_),
    .C1(_06547_),
    .C2(_06407_),
    .ZN(_06640_));
 OAI21_X1 _30151_ (.A(_06496_),
    .B1(_06474_),
    .B2(_06533_),
    .ZN(_06641_));
 NAND3_X1 _30152_ (.A1(_06464_),
    .A2(_06468_),
    .A3(_06641_),
    .ZN(_06642_));
 NOR4_X2 _30153_ (.A1(_06505_),
    .A2(_06588_),
    .A3(_06590_),
    .A4(_06596_),
    .ZN(_06643_));
 NOR2_X1 _30154_ (.A1(_22546_),
    .A2(_19434_),
    .ZN(_06644_));
 OR3_X1 _30155_ (.A1(_06642_),
    .A2(_06643_),
    .A3(_06644_),
    .ZN(_06645_));
 AND3_X1 _30156_ (.A1(_06636_),
    .A2(_06640_),
    .A3(_06645_),
    .ZN(_06646_));
 MUX2_X1 _30157_ (.A(_06298_),
    .B(_06352_),
    .S(_06420_),
    .Z(_06647_));
 NOR2_X1 _30158_ (.A1(_06464_),
    .A2(_06647_),
    .ZN(_06648_));
 OAI21_X1 _30159_ (.A(_06456_),
    .B1(_06298_),
    .B2(_06420_),
    .ZN(_06649_));
 AOI221_X4 _30160_ (.A(_06648_),
    .B1(_06649_),
    .B2(_06643_),
    .C1(_06644_),
    .C2(_06464_),
    .ZN(_06650_));
 MUX2_X1 _30161_ (.A(_06391_),
    .B(_06353_),
    .S(_06421_),
    .Z(_06651_));
 OAI33_X1 _30162_ (.A1(_06505_),
    .A2(_06599_),
    .A3(_06625_),
    .B1(_06651_),
    .B2(_06480_),
    .B3(_06464_),
    .ZN(_06652_));
 AND2_X1 _30163_ (.A1(_06465_),
    .A2(_06652_),
    .ZN(_06653_));
 AOI21_X1 _30164_ (.A(_06578_),
    .B1(_06460_),
    .B2(_06459_),
    .ZN(_06654_));
 MUX2_X1 _30165_ (.A(_06349_),
    .B(_06392_),
    .S(_06421_),
    .Z(_06655_));
 MUX2_X1 _30166_ (.A(_06654_),
    .B(_06655_),
    .S(_06456_),
    .Z(_06656_));
 OR3_X1 _30167_ (.A1(_06478_),
    .A2(_06555_),
    .A3(_06560_),
    .ZN(_06657_));
 OAI33_X1 _30168_ (.A1(_14204_),
    .A2(_06386_),
    .A3(_06457_),
    .B1(_06454_),
    .B2(_06312_),
    .B3(_06330_),
    .ZN(_06658_));
 AND4_X1 _30169_ (.A1(_06538_),
    .A2(_06442_),
    .A3(_06444_),
    .A4(_06445_),
    .ZN(_06659_));
 AOI21_X1 _30170_ (.A(_06658_),
    .B1(_06659_),
    .B2(_06554_),
    .ZN(_06660_));
 MUX2_X1 _30171_ (.A(_06293_),
    .B(_06409_),
    .S(_06420_),
    .Z(_06661_));
 AOI22_X2 _30172_ (.A1(_06660_),
    .A2(_06598_),
    .B1(_06661_),
    .B2(_06456_),
    .ZN(_06662_));
 INV_X1 _30173_ (.A(_06579_),
    .ZN(_06663_));
 AOI221_X2 _30174_ (.A(_06656_),
    .B1(_06657_),
    .B2(_06662_),
    .C1(_06544_),
    .C2(_06663_),
    .ZN(_06664_));
 MUX2_X1 _30175_ (.A(_06290_),
    .B(_06348_),
    .S(_06547_),
    .Z(_06665_));
 MUX2_X1 _30176_ (.A(_06610_),
    .B(_06535_),
    .S(_06402_),
    .Z(_06666_));
 NAND2_X1 _30177_ (.A1(_06525_),
    .A2(_06504_),
    .ZN(_06667_));
 NAND2_X1 _30178_ (.A1(_14204_),
    .A2(_06504_),
    .ZN(_06668_));
 NAND2_X1 _30179_ (.A1(_06507_),
    .A2(_06460_),
    .ZN(_06669_));
 MUX2_X1 _30180_ (.A(_06543_),
    .B(_06669_),
    .S(_06402_),
    .Z(_06670_));
 OAI222_X4 _30181_ (.A1(_06464_),
    .A2(_06665_),
    .B1(_06666_),
    .B2(_06667_),
    .C1(_06668_),
    .C2(_06670_),
    .ZN(_06671_));
 NAND4_X2 _30182_ (.A1(_06650_),
    .A2(_06653_),
    .A3(_06664_),
    .A4(_06671_),
    .ZN(_06672_));
 NOR3_X1 _30183_ (.A1(_06634_),
    .A2(_06646_),
    .A3(_06672_),
    .ZN(_06673_));
 XNOR2_X2 _30184_ (.A(_06549_),
    .B(_06673_),
    .ZN(_22556_));
 MUX2_X1 _30185_ (.A(_06503_),
    .B(_22553_),
    .S(_22556_),
    .Z(_06674_));
 NAND2_X1 _30186_ (.A1(_06486_),
    .A2(_06674_),
    .ZN(_06675_));
 AOI21_X1 _30187_ (.A(_06482_),
    .B1(_06484_),
    .B2(_06675_),
    .ZN(_00176_));
 NOR2_X1 _30188_ (.A1(\g_reduce0[14].adder.x[1] ),
    .A2(_06481_),
    .ZN(_06676_));
 AOI21_X1 _30189_ (.A(_06483_),
    .B1(_06064_),
    .B2(\g_reduce0[12].adder.x[1] ),
    .ZN(_06677_));
 OR2_X1 _30190_ (.A1(_22553_),
    .A2(_22556_),
    .ZN(_06678_));
 AND2_X1 _30191_ (.A1(_06642_),
    .A2(_06650_),
    .ZN(_06679_));
 XNOR2_X1 _30192_ (.A(_22552_),
    .B(_06679_),
    .ZN(_06680_));
 NAND2_X1 _30193_ (.A1(_22556_),
    .A2(_06680_),
    .ZN(_06681_));
 NAND3_X1 _30194_ (.A1(_06486_),
    .A2(_06678_),
    .A3(_06681_),
    .ZN(_06682_));
 AOI21_X1 _30195_ (.A(_06676_),
    .B1(_06677_),
    .B2(_06682_),
    .ZN(_00183_));
 OAI21_X1 _30196_ (.A(_06061_),
    .B1(_06486_),
    .B2(\g_reduce0[12].adder.x[2] ),
    .ZN(_06683_));
 AND2_X1 _30197_ (.A1(_06650_),
    .A2(_06653_),
    .ZN(_06684_));
 AOI21_X1 _30198_ (.A(_06656_),
    .B1(_06663_),
    .B2(_06544_),
    .ZN(_06685_));
 XOR2_X1 _30199_ (.A(_06684_),
    .B(_06685_),
    .Z(_06686_));
 NAND2_X1 _30200_ (.A1(_06642_),
    .A2(_06686_),
    .ZN(_06687_));
 MUX2_X1 _30201_ (.A(_06680_),
    .B(_06687_),
    .S(_22556_),
    .Z(_06688_));
 AOI21_X1 _30202_ (.A(_06683_),
    .B1(_06688_),
    .B2(_06486_),
    .ZN(_06689_));
 AOI21_X1 _30203_ (.A(_06689_),
    .B1(_06483_),
    .B2(\g_reduce0[14].adder.x[2] ),
    .ZN(_06690_));
 INV_X1 _30204_ (.A(_06690_),
    .ZN(_00184_));
 OAI21_X1 _30205_ (.A(_06061_),
    .B1(_06486_),
    .B2(\g_reduce0[12].adder.x[3] ),
    .ZN(_06691_));
 NAND2_X1 _30206_ (.A1(_06662_),
    .A2(_06657_),
    .ZN(_06692_));
 NAND3_X1 _30207_ (.A1(_22552_),
    .A2(_06685_),
    .A3(_06679_),
    .ZN(_06693_));
 XOR2_X1 _30208_ (.A(_06692_),
    .B(_06693_),
    .Z(_06694_));
 MUX2_X1 _30209_ (.A(_06687_),
    .B(_06694_),
    .S(_22556_),
    .Z(_06695_));
 AOI21_X1 _30210_ (.A(_06691_),
    .B1(_06695_),
    .B2(_06486_),
    .ZN(_06696_));
 AOI21_X1 _30211_ (.A(_06696_),
    .B1(_06483_),
    .B2(\g_reduce0[14].adder.x[3] ),
    .ZN(_06697_));
 INV_X1 _30212_ (.A(_06697_),
    .ZN(_00185_));
 NOR2_X4 _30213_ (.A1(_06483_),
    .A2(_06486_),
    .ZN(_06698_));
 AOI22_X2 _30214_ (.A1(\g_reduce0[14].adder.x[4] ),
    .A2(_06483_),
    .B1(_06698_),
    .B2(\g_reduce0[12].adder.x[4] ),
    .ZN(_06699_));
 NAND2_X1 _30215_ (.A1(_06684_),
    .A2(_06664_),
    .ZN(_06700_));
 XOR2_X1 _30216_ (.A(_06700_),
    .B(_06671_),
    .Z(_06701_));
 MUX2_X1 _30217_ (.A(_06694_),
    .B(_06701_),
    .S(_22556_),
    .Z(_06702_));
 NAND2_X1 _30218_ (.A1(_06061_),
    .A2(_06485_),
    .ZN(_06703_));
 OAI21_X1 _30219_ (.A(_06699_),
    .B1(_06702_),
    .B2(_06703_),
    .ZN(_00186_));
 INV_X1 _30220_ (.A(_06703_),
    .ZN(_06704_));
 INV_X1 _30221_ (.A(_06549_),
    .ZN(_06705_));
 OAI21_X1 _30222_ (.A(_06704_),
    .B1(_06701_),
    .B2(_06705_),
    .ZN(_06706_));
 NAND4_X2 _30223_ (.A1(_22552_),
    .A2(_06664_),
    .A3(_06671_),
    .A4(_06679_),
    .ZN(_06707_));
 XNOR2_X1 _30224_ (.A(_06609_),
    .B(_06707_),
    .ZN(_06708_));
 AOI21_X1 _30225_ (.A(_06706_),
    .B1(_06708_),
    .B2(_22556_),
    .ZN(_06709_));
 NAND2_X1 _30226_ (.A1(_06061_),
    .A2(_06064_),
    .ZN(_06710_));
 OAI22_X2 _30227_ (.A1(\g_reduce0[14].adder.x[5] ),
    .A2(_06481_),
    .B1(_06710_),
    .B2(\g_reduce0[12].adder.x[5] ),
    .ZN(_06711_));
 NOR2_X1 _30228_ (.A1(_06709_),
    .A2(_06711_),
    .ZN(_00187_));
 INV_X1 _30229_ (.A(_06708_),
    .ZN(_06712_));
 NAND4_X1 _30230_ (.A1(_06609_),
    .A2(_06684_),
    .A3(_06664_),
    .A4(_06671_),
    .ZN(_06713_));
 XOR2_X1 _30231_ (.A(_06582_),
    .B(_06713_),
    .Z(_06714_));
 OAI221_X1 _30232_ (.A(_06704_),
    .B1(_06712_),
    .B2(_22556_),
    .C1(_06714_),
    .C2(_06549_),
    .ZN(_06715_));
 OAI22_X1 _30233_ (.A1(\g_reduce0[14].adder.x[6] ),
    .A2(_06481_),
    .B1(_06710_),
    .B2(\g_reduce0[12].adder.x[6] ),
    .ZN(_06716_));
 INV_X1 _30234_ (.A(_06716_),
    .ZN(_06717_));
 AND2_X1 _30235_ (.A1(_06715_),
    .A2(_06717_),
    .ZN(_00188_));
 AOI22_X4 _30236_ (.A1(\g_reduce0[14].adder.x[7] ),
    .A2(_06483_),
    .B1(_06698_),
    .B2(\g_reduce0[12].adder.x[7] ),
    .ZN(_06718_));
 NAND2_X1 _30237_ (.A1(_06582_),
    .A2(_06609_),
    .ZN(_06719_));
 NOR2_X1 _30238_ (.A1(_06719_),
    .A2(_06707_),
    .ZN(_06720_));
 XNOR2_X1 _30239_ (.A(_06577_),
    .B(_06720_),
    .ZN(_06721_));
 MUX2_X1 _30240_ (.A(_06714_),
    .B(_06721_),
    .S(_22556_),
    .Z(_06722_));
 OAI21_X1 _30241_ (.A(_06718_),
    .B1(_06722_),
    .B2(_06703_),
    .ZN(_00189_));
 OAI21_X1 _30242_ (.A(_06549_),
    .B1(_06673_),
    .B2(_06721_),
    .ZN(_06723_));
 NAND3_X1 _30243_ (.A1(_06577_),
    .A2(_06582_),
    .A3(_06609_),
    .ZN(_06724_));
 NOR2_X1 _30244_ (.A1(_06724_),
    .A2(_06672_),
    .ZN(_06725_));
 OR3_X1 _30245_ (.A1(_06549_),
    .A2(_06633_),
    .A3(_06725_),
    .ZN(_06726_));
 INV_X1 _30246_ (.A(_06646_),
    .ZN(_06727_));
 OAI21_X1 _30247_ (.A(_06707_),
    .B1(_06727_),
    .B2(_06549_),
    .ZN(_06728_));
 NAND2_X1 _30248_ (.A1(_06633_),
    .A2(_06671_),
    .ZN(_06729_));
 NOR3_X1 _30249_ (.A1(_06724_),
    .A2(_06700_),
    .A3(_06729_),
    .ZN(_06730_));
 AOI21_X1 _30250_ (.A(_06703_),
    .B1(_06728_),
    .B2(_06730_),
    .ZN(_06731_));
 NAND3_X1 _30251_ (.A1(_06723_),
    .A2(_06726_),
    .A3(_06731_),
    .ZN(_06732_));
 AOI22_X4 _30252_ (.A1(\g_reduce0[14].adder.x[8] ),
    .A2(_06483_),
    .B1(_06698_),
    .B2(\g_reduce0[12].adder.x[8] ),
    .ZN(_06733_));
 NAND2_X1 _30253_ (.A1(_06732_),
    .A2(_06733_),
    .ZN(_00190_));
 NAND2_X1 _30254_ (.A1(\g_reduce0[14].adder.x[9] ),
    .A2(_06483_),
    .ZN(_06734_));
 OAI21_X1 _30255_ (.A(_06481_),
    .B1(_06486_),
    .B2(\g_reduce0[12].adder.x[9] ),
    .ZN(_06735_));
 XNOR2_X1 _30256_ (.A(_06633_),
    .B(_06725_),
    .ZN(_06736_));
 OAI21_X1 _30257_ (.A(_06485_),
    .B1(_06705_),
    .B2(_06736_),
    .ZN(_06737_));
 NOR2_X1 _30258_ (.A1(_06634_),
    .A2(_06707_),
    .ZN(_06738_));
 NOR2_X1 _30259_ (.A1(_06646_),
    .A2(_06738_),
    .ZN(_06739_));
 NOR2_X1 _30260_ (.A1(_06634_),
    .A2(_06672_),
    .ZN(_06740_));
 XNOR2_X1 _30261_ (.A(_06549_),
    .B(_06740_),
    .ZN(_06741_));
 NOR2_X1 _30262_ (.A1(_06549_),
    .A2(_06727_),
    .ZN(_06742_));
 AOI221_X2 _30263_ (.A(_06737_),
    .B1(_06739_),
    .B2(_06741_),
    .C1(_06742_),
    .C2(_06738_),
    .ZN(_06743_));
 OAI21_X1 _30264_ (.A(_06734_),
    .B1(_06735_),
    .B2(_06743_),
    .ZN(_00191_));
 MUX2_X1 _30265_ (.A(\g_reduce0[12].adder.x[10] ),
    .B(_22558_),
    .S(_06486_),
    .Z(_06744_));
 MUX2_X1 _30266_ (.A(\g_reduce0[14].adder.x[10] ),
    .B(_06744_),
    .S(_06481_),
    .Z(_00177_));
 MUX2_X1 _30267_ (.A(_06057_),
    .B(_19432_),
    .S(_06486_),
    .Z(_06745_));
 MUX2_X1 _30268_ (.A(\g_reduce0[14].adder.x[11] ),
    .B(_06745_),
    .S(_06481_),
    .Z(_00178_));
 XNOR2_X1 _30269_ (.A(_14207_),
    .B(_19436_),
    .ZN(_06746_));
 MUX2_X2 _30270_ (.A(_22432_),
    .B(_00612_),
    .S(_06102_),
    .Z(_06747_));
 NAND2_X1 _30271_ (.A1(_06420_),
    .A2(_19425_),
    .ZN(_06748_));
 XOR2_X1 _30272_ (.A(_06747_),
    .B(_06748_),
    .Z(_06749_));
 MUX2_X1 _30273_ (.A(_06746_),
    .B(_06749_),
    .S(_06456_),
    .Z(_06750_));
 XOR2_X1 _30274_ (.A(_19431_),
    .B(_06750_),
    .Z(_06751_));
 MUX2_X1 _30275_ (.A(_06058_),
    .B(_06751_),
    .S(_06485_),
    .Z(_06752_));
 MUX2_X1 _30276_ (.A(\g_reduce0[14].adder.x[12] ),
    .B(_06752_),
    .S(_06481_),
    .Z(_00179_));
 INV_X1 _30277_ (.A(_19435_),
    .ZN(_06753_));
 INV_X1 _30278_ (.A(_14206_),
    .ZN(_06754_));
 AOI21_X1 _30279_ (.A(_19427_),
    .B1(_19428_),
    .B2(_06754_),
    .ZN(_06755_));
 INV_X1 _30280_ (.A(_19436_),
    .ZN(_06756_));
 OAI21_X1 _30281_ (.A(_06753_),
    .B1(_06755_),
    .B2(_06756_),
    .ZN(_06757_));
 XOR2_X1 _30282_ (.A(_19440_),
    .B(_06757_),
    .Z(_06758_));
 MUX2_X1 _30283_ (.A(_22429_),
    .B(_00615_),
    .S(_06102_),
    .Z(_06759_));
 NOR4_X1 _30284_ (.A1(_06547_),
    .A2(_22554_),
    .A3(_14205_),
    .A4(_06747_),
    .ZN(_06760_));
 XNOR2_X1 _30285_ (.A(_06759_),
    .B(_06760_),
    .ZN(_06761_));
 MUX2_X1 _30286_ (.A(_06758_),
    .B(_06761_),
    .S(_06456_),
    .Z(_06762_));
 NOR2_X1 _30287_ (.A1(_06547_),
    .A2(_19426_),
    .ZN(_06763_));
 AOI21_X1 _30288_ (.A(_06763_),
    .B1(_14205_),
    .B2(_06547_),
    .ZN(_06764_));
 NOR2_X1 _30289_ (.A1(_06499_),
    .A2(_06764_),
    .ZN(_06765_));
 AOI21_X2 _30290_ (.A(_06765_),
    .B1(_06499_),
    .B2(_14208_),
    .ZN(_19430_));
 NAND3_X1 _30291_ (.A1(_19429_),
    .A2(_06750_),
    .A3(_19430_),
    .ZN(_06766_));
 XNOR2_X1 _30292_ (.A(_06762_),
    .B(_06766_),
    .ZN(_06767_));
 MUX2_X1 _30293_ (.A(\g_reduce0[12].adder.x[13] ),
    .B(_06767_),
    .S(_06485_),
    .Z(_06768_));
 MUX2_X1 _30294_ (.A(\g_reduce0[14].adder.x[13] ),
    .B(_06768_),
    .S(_06481_),
    .Z(_00180_));
 INV_X1 _30295_ (.A(_22430_),
    .ZN(_06769_));
 AOI22_X1 _30296_ (.A1(_06069_),
    .A2(_22433_),
    .B1(_06071_),
    .B2(_06068_),
    .ZN(_06770_));
 AOI21_X1 _30297_ (.A(_06073_),
    .B1(_06769_),
    .B2(_06770_),
    .ZN(_06771_));
 NOR2_X1 _30298_ (.A1(_22475_),
    .A2(_06771_),
    .ZN(_06772_));
 INV_X1 _30299_ (.A(_06772_),
    .ZN(_06773_));
 OR2_X1 _30300_ (.A1(_06062_),
    .A2(_06773_),
    .ZN(_06774_));
 NAND2_X1 _30301_ (.A1(_06059_),
    .A2(_06774_),
    .ZN(_06775_));
 NOR4_X1 _30302_ (.A1(_06499_),
    .A2(_06747_),
    .A3(_06748_),
    .A4(_06759_),
    .ZN(_06776_));
 OAI21_X1 _30303_ (.A(_06753_),
    .B1(_06756_),
    .B2(_14207_),
    .ZN(_06777_));
 AOI21_X1 _30304_ (.A(_19439_),
    .B1(_06777_),
    .B2(_19440_),
    .ZN(_06778_));
 AOI21_X1 _30305_ (.A(_06776_),
    .B1(_06778_),
    .B2(_06499_),
    .ZN(_06779_));
 NAND3_X1 _30306_ (.A1(_19431_),
    .A2(_06750_),
    .A3(_06762_),
    .ZN(_06780_));
 XNOR2_X2 _30307_ (.A(_06779_),
    .B(_06780_),
    .ZN(_06781_));
 MUX2_X1 _30308_ (.A(_06775_),
    .B(_06774_),
    .S(_06781_),
    .Z(_06782_));
 OAI22_X1 _30309_ (.A1(_06062_),
    .A2(_06481_),
    .B1(_06064_),
    .B2(_06782_),
    .ZN(_06783_));
 NOR2_X1 _30310_ (.A1(_06059_),
    .A2(_06483_),
    .ZN(_06784_));
 AOI21_X1 _30311_ (.A(_06064_),
    .B1(_06773_),
    .B2(_06781_),
    .ZN(_06785_));
 NAND2_X1 _30312_ (.A1(_06062_),
    .A2(_06772_),
    .ZN(_06786_));
 OAI21_X1 _30313_ (.A(_06785_),
    .B1(_06786_),
    .B2(_06781_),
    .ZN(_06787_));
 AOI21_X1 _30314_ (.A(_06783_),
    .B1(_06784_),
    .B2(_06787_),
    .ZN(_00181_));
 CLKBUF_X2 _30315_ (.A(_19464_),
    .Z(_06788_));
 AOI21_X1 _30316_ (.A(_19463_),
    .B1(_06788_),
    .B2(_19465_),
    .ZN(_06789_));
 BUF_X1 _30317_ (.A(_19466_),
    .Z(_06790_));
 NAND2_X1 _30318_ (.A1(_06788_),
    .A2(_06790_),
    .ZN(_06791_));
 CLKBUF_X2 _30319_ (.A(_19469_),
    .Z(_06792_));
 AOI21_X1 _30320_ (.A(_19467_),
    .B1(_19468_),
    .B2(_06792_),
    .ZN(_06793_));
 OAI21_X1 _30321_ (.A(_06789_),
    .B1(_06791_),
    .B2(_06793_),
    .ZN(_06794_));
 INV_X1 _30322_ (.A(_19471_),
    .ZN(_06795_));
 CLKBUF_X2 _30323_ (.A(_19473_),
    .Z(_06796_));
 INV_X1 _30324_ (.A(_19475_),
    .ZN(_06797_));
 AOI21_X1 _30325_ (.A(_19477_),
    .B1(_19478_),
    .B2(_19479_),
    .ZN(_06798_));
 INV_X1 _30326_ (.A(_19476_),
    .ZN(_06799_));
 OAI21_X1 _30327_ (.A(_06797_),
    .B1(_06798_),
    .B2(_06799_),
    .ZN(_06800_));
 CLKBUF_X2 _30328_ (.A(_19474_),
    .Z(_06801_));
 AOI21_X1 _30329_ (.A(_06796_),
    .B1(_06800_),
    .B2(_06801_),
    .ZN(_06802_));
 INV_X1 _30330_ (.A(_19472_),
    .ZN(_06803_));
 OAI21_X2 _30331_ (.A(_06795_),
    .B1(_06802_),
    .B2(_06803_),
    .ZN(_06804_));
 INV_X1 _30332_ (.A(_19468_),
    .ZN(_06805_));
 CLKBUF_X2 _30333_ (.A(_19470_),
    .Z(_06806_));
 INV_X1 _30334_ (.A(_06806_),
    .ZN(_06807_));
 NOR3_X2 _30335_ (.A1(_06805_),
    .A2(_06807_),
    .A3(_06791_),
    .ZN(_06808_));
 AOI21_X2 _30336_ (.A(_06794_),
    .B1(_06804_),
    .B2(_06808_),
    .ZN(_06809_));
 XNOR2_X2 _30337_ (.A(_19462_),
    .B(_06809_),
    .ZN(_06810_));
 INV_X1 _30338_ (.A(_06810_),
    .ZN(_06811_));
 INV_X1 _30339_ (.A(_19467_),
    .ZN(_06812_));
 AOI21_X1 _30340_ (.A(_06792_),
    .B1(_06806_),
    .B2(_06804_),
    .ZN(_06813_));
 OAI21_X2 _30341_ (.A(_06812_),
    .B1(_06813_),
    .B2(_06805_),
    .ZN(_06814_));
 XNOR2_X1 _30342_ (.A(_06790_),
    .B(_06814_),
    .ZN(_06815_));
 XNOR2_X1 _30343_ (.A(_06807_),
    .B(_06804_),
    .ZN(_06816_));
 INV_X1 _30344_ (.A(_19461_),
    .ZN(_06817_));
 INV_X1 _30345_ (.A(_19462_),
    .ZN(_06818_));
 AOI21_X1 _30346_ (.A(_19465_),
    .B1(_06790_),
    .B2(_19467_),
    .ZN(_06819_));
 INV_X1 _30347_ (.A(_06819_),
    .ZN(_06820_));
 AOI21_X1 _30348_ (.A(_19463_),
    .B1(_06820_),
    .B2(_06788_),
    .ZN(_06821_));
 OAI21_X1 _30349_ (.A(_06817_),
    .B1(_06818_),
    .B2(_06821_),
    .ZN(_06822_));
 INV_X1 _30350_ (.A(_06788_),
    .ZN(_06823_));
 NAND2_X1 _30351_ (.A1(_06790_),
    .A2(_19468_),
    .ZN(_06824_));
 NOR3_X2 _30352_ (.A1(_06818_),
    .A2(_06823_),
    .A3(_06824_),
    .ZN(_06825_));
 AOI21_X2 _30353_ (.A(_06792_),
    .B1(_06806_),
    .B2(_19471_),
    .ZN(_06826_));
 OAI21_X1 _30354_ (.A(_06797_),
    .B1(_06799_),
    .B2(_14214_),
    .ZN(_06827_));
 AOI21_X1 _30355_ (.A(_06796_),
    .B1(_06827_),
    .B2(_06801_),
    .ZN(_06828_));
 NAND2_X1 _30356_ (.A1(_06806_),
    .A2(_19472_),
    .ZN(_06829_));
 NOR2_X1 _30357_ (.A1(_06828_),
    .A2(_06829_),
    .ZN(_06830_));
 INV_X1 _30358_ (.A(_06830_),
    .ZN(_06831_));
 NAND2_X1 _30359_ (.A1(_06826_),
    .A2(_06831_),
    .ZN(_06832_));
 AOI21_X1 _30360_ (.A(_06822_),
    .B1(_06825_),
    .B2(_06832_),
    .ZN(_06833_));
 XNOR2_X1 _30361_ (.A(_19460_),
    .B(_06833_),
    .ZN(_19494_));
 XNOR2_X1 _30362_ (.A(_06803_),
    .B(_06828_),
    .ZN(_06834_));
 XNOR2_X1 _30363_ (.A(_06801_),
    .B(_06800_),
    .ZN(_06835_));
 AOI21_X1 _30364_ (.A(_06807_),
    .B1(_06803_),
    .B2(_06795_),
    .ZN(_06836_));
 NOR2_X1 _30365_ (.A1(_06792_),
    .A2(_06836_),
    .ZN(_06837_));
 XNOR2_X1 _30366_ (.A(_06805_),
    .B(_06837_),
    .ZN(_06838_));
 XNOR2_X1 _30367_ (.A(_14214_),
    .B(_19476_),
    .ZN(_06839_));
 NOR4_X1 _30368_ (.A1(_14215_),
    .A2(\g_row[0].g_col[0].mult.adder.a[0] ),
    .A3(_19480_),
    .A4(_06839_),
    .ZN(_06840_));
 NAND4_X1 _30369_ (.A1(_06834_),
    .A2(_06835_),
    .A3(_06838_),
    .A4(_06840_),
    .ZN(_06841_));
 OAI21_X1 _30370_ (.A(_06819_),
    .B1(_06824_),
    .B2(_06826_),
    .ZN(_06842_));
 NOR2_X1 _30371_ (.A1(_06824_),
    .A2(_06831_),
    .ZN(_06843_));
 NOR2_X1 _30372_ (.A1(_06842_),
    .A2(_06843_),
    .ZN(_06844_));
 XNOR2_X1 _30373_ (.A(_06788_),
    .B(_06844_),
    .ZN(_06845_));
 NOR4_X1 _30374_ (.A1(_06816_),
    .A2(_19494_),
    .A3(_06841_),
    .A4(_06845_),
    .ZN(_06846_));
 AND2_X1 _30375_ (.A1(_06815_),
    .A2(_06846_),
    .ZN(_06847_));
 NOR2_X1 _30376_ (.A1(_06811_),
    .A2(_06847_),
    .ZN(_19495_));
 INV_X1 _30377_ (.A(_19441_),
    .ZN(_06848_));
 INV_X1 _30378_ (.A(_19442_),
    .ZN(_06849_));
 INV_X1 _30379_ (.A(_19445_),
    .ZN(_06850_));
 INV_X1 _30380_ (.A(_19446_),
    .ZN(_06851_));
 INV_X1 _30381_ (.A(_19451_),
    .ZN(_06852_));
 BUF_X2 _30382_ (.A(_19454_),
    .Z(_06853_));
 AOI21_X2 _30383_ (.A(_19453_),
    .B1(_06853_),
    .B2(_19455_),
    .ZN(_06854_));
 BUF_X2 _30384_ (.A(_19452_),
    .Z(_06855_));
 INV_X1 _30385_ (.A(_06855_),
    .ZN(_06856_));
 OAI21_X1 _30386_ (.A(_06852_),
    .B1(_06854_),
    .B2(_06856_),
    .ZN(_06857_));
 AOI21_X2 _30387_ (.A(_19449_),
    .B1(_19450_),
    .B2(_06857_),
    .ZN(_06858_));
 BUF_X2 _30388_ (.A(_19458_),
    .Z(_06859_));
 AND2_X1 _30389_ (.A1(_06859_),
    .A2(_19460_),
    .ZN(_06860_));
 AOI21_X1 _30390_ (.A(_19463_),
    .B1(_06842_),
    .B2(_06788_),
    .ZN(_06861_));
 OAI21_X1 _30391_ (.A(_06817_),
    .B1(_06818_),
    .B2(_06861_),
    .ZN(_06862_));
 AOI221_X2 _30392_ (.A(_19457_),
    .B1(_06859_),
    .B2(_19459_),
    .C1(_06860_),
    .C2(_06862_),
    .ZN(_06863_));
 BUF_X2 _30393_ (.A(_19456_),
    .Z(_06864_));
 NAND4_X2 _30394_ (.A1(_19450_),
    .A2(_06855_),
    .A3(_06853_),
    .A4(_06864_),
    .ZN(_06865_));
 OAI21_X1 _30395_ (.A(_06858_),
    .B1(_06863_),
    .B2(_06865_),
    .ZN(_06866_));
 BUF_X2 _30396_ (.A(_19448_),
    .Z(_06867_));
 AOI21_X1 _30397_ (.A(_19447_),
    .B1(_06866_),
    .B2(_06867_),
    .ZN(_06868_));
 OAI21_X1 _30398_ (.A(_06850_),
    .B1(_06851_),
    .B2(_06868_),
    .ZN(_06869_));
 AOI21_X2 _30399_ (.A(_19443_),
    .B1(_19444_),
    .B2(_06869_),
    .ZN(_06870_));
 OAI21_X4 _30400_ (.A(_06848_),
    .B1(_06849_),
    .B2(_06870_),
    .ZN(_06871_));
 INV_X1 _30401_ (.A(_19453_),
    .ZN(_06872_));
 INV_X1 _30402_ (.A(_06853_),
    .ZN(_06873_));
 AOI21_X1 _30403_ (.A(_19455_),
    .B1(_06864_),
    .B2(_19457_),
    .ZN(_06874_));
 OAI21_X1 _30404_ (.A(_06872_),
    .B1(_06873_),
    .B2(_06874_),
    .ZN(_06875_));
 AOI21_X1 _30405_ (.A(_19451_),
    .B1(_06875_),
    .B2(_06855_),
    .ZN(_06876_));
 NAND4_X1 _30406_ (.A1(_06855_),
    .A2(_06853_),
    .A3(_06864_),
    .A4(_06859_),
    .ZN(_06877_));
 AOI21_X1 _30407_ (.A(_19459_),
    .B1(_19460_),
    .B2(_19461_),
    .ZN(_06878_));
 NAND2_X1 _30408_ (.A1(_19460_),
    .A2(_19462_),
    .ZN(_06879_));
 OAI21_X1 _30409_ (.A(_06878_),
    .B1(_06879_),
    .B2(_06789_),
    .ZN(_06880_));
 NOR2_X1 _30410_ (.A1(_06791_),
    .A2(_06879_),
    .ZN(_06881_));
 INV_X1 _30411_ (.A(_06796_),
    .ZN(_06882_));
 OAI21_X1 _30412_ (.A(_06795_),
    .B1(_06882_),
    .B2(_06803_),
    .ZN(_06883_));
 AOI21_X1 _30413_ (.A(_06792_),
    .B1(_06806_),
    .B2(_06883_),
    .ZN(_06884_));
 OAI21_X1 _30414_ (.A(_06812_),
    .B1(_06884_),
    .B2(_06805_),
    .ZN(_06885_));
 AOI21_X1 _30415_ (.A(_06880_),
    .B1(_06881_),
    .B2(_06885_),
    .ZN(_06886_));
 OAI21_X1 _30416_ (.A(_06876_),
    .B1(_06877_),
    .B2(_06886_),
    .ZN(_06887_));
 AOI21_X1 _30417_ (.A(_19449_),
    .B1(_19450_),
    .B2(_06887_),
    .ZN(_06888_));
 INV_X1 _30418_ (.A(_06888_),
    .ZN(_06889_));
 AOI21_X1 _30419_ (.A(_19447_),
    .B1(_06889_),
    .B2(_06867_),
    .ZN(_06890_));
 OAI21_X1 _30420_ (.A(_06850_),
    .B1(_06851_),
    .B2(_06890_),
    .ZN(_06891_));
 AOI21_X1 _30421_ (.A(_19443_),
    .B1(_19444_),
    .B2(_06891_),
    .ZN(_06892_));
 XNOR2_X1 _30422_ (.A(_19442_),
    .B(_06892_),
    .ZN(_06893_));
 NAND2_X1 _30423_ (.A1(_06825_),
    .A2(_06860_),
    .ZN(_06894_));
 OAI21_X2 _30424_ (.A(_06863_),
    .B1(_06894_),
    .B2(_06831_),
    .ZN(_06895_));
 INV_X1 _30425_ (.A(_06895_),
    .ZN(_06896_));
 OAI21_X2 _30426_ (.A(_06858_),
    .B1(_06865_),
    .B2(_06896_),
    .ZN(_06897_));
 XOR2_X2 _30427_ (.A(_06867_),
    .B(_06897_),
    .Z(_06898_));
 INV_X1 _30428_ (.A(_19449_),
    .ZN(_06899_));
 INV_X1 _30429_ (.A(_19450_),
    .ZN(_06900_));
 NAND2_X1 _30430_ (.A1(_06864_),
    .A2(_06859_),
    .ZN(_06901_));
 OAI21_X1 _30431_ (.A(_06874_),
    .B1(_06901_),
    .B2(_06878_),
    .ZN(_06902_));
 INV_X1 _30432_ (.A(_19477_),
    .ZN(_06903_));
 OAI21_X1 _30433_ (.A(_06797_),
    .B1(_06903_),
    .B2(_06799_),
    .ZN(_06904_));
 AOI21_X1 _30434_ (.A(_06796_),
    .B1(_06904_),
    .B2(_06801_),
    .ZN(_06905_));
 OAI21_X1 _30435_ (.A(_06795_),
    .B1(_06905_),
    .B2(_06803_),
    .ZN(_06906_));
 AOI21_X1 _30436_ (.A(_06794_),
    .B1(_06808_),
    .B2(_06906_),
    .ZN(_06907_));
 NOR3_X1 _30437_ (.A1(_06901_),
    .A2(_06879_),
    .A3(_06907_),
    .ZN(_06908_));
 OAI21_X1 _30438_ (.A(_06853_),
    .B1(_06902_),
    .B2(_06908_),
    .ZN(_06909_));
 NAND2_X1 _30439_ (.A1(_06872_),
    .A2(_06909_),
    .ZN(_06910_));
 AOI21_X1 _30440_ (.A(_19451_),
    .B1(_06910_),
    .B2(_06855_),
    .ZN(_06911_));
 OAI21_X1 _30441_ (.A(_06899_),
    .B1(_06900_),
    .B2(_06911_),
    .ZN(_06912_));
 AOI21_X2 _30442_ (.A(_19447_),
    .B1(_06912_),
    .B2(_06867_),
    .ZN(_06913_));
 XNOR2_X2 _30443_ (.A(_19446_),
    .B(_06913_),
    .ZN(_06914_));
 AOI21_X2 _30444_ (.A(_19457_),
    .B1(_06859_),
    .B2(_19459_),
    .ZN(_06915_));
 NAND2_X1 _30445_ (.A1(_06853_),
    .A2(_06864_),
    .ZN(_06916_));
 NAND3_X1 _30446_ (.A1(_06853_),
    .A2(_06864_),
    .A3(_06860_),
    .ZN(_06917_));
 OAI221_X2 _30447_ (.A(_06854_),
    .B1(_06915_),
    .B2(_06916_),
    .C1(_06917_),
    .C2(_06833_),
    .ZN(_06918_));
 XNOR2_X2 _30448_ (.A(_06856_),
    .B(_06918_),
    .ZN(_06919_));
 AOI21_X2 _30449_ (.A(_06880_),
    .B1(_06881_),
    .B2(_06814_),
    .ZN(_06920_));
 XNOR2_X2 _30450_ (.A(_06859_),
    .B(_06920_),
    .ZN(_06921_));
 AND3_X1 _30451_ (.A1(_06810_),
    .A2(_19494_),
    .A3(_06921_),
    .ZN(_06922_));
 NOR3_X1 _30452_ (.A1(_06809_),
    .A2(_06901_),
    .A3(_06879_),
    .ZN(_06923_));
 NOR2_X1 _30453_ (.A1(_06902_),
    .A2(_06923_),
    .ZN(_06924_));
 XNOR2_X2 _30454_ (.A(_06873_),
    .B(_06924_),
    .ZN(_06925_));
 INV_X1 _30455_ (.A(_06925_),
    .ZN(_06926_));
 XOR2_X2 _30456_ (.A(_06864_),
    .B(_06895_),
    .Z(_06927_));
 AND3_X1 _30457_ (.A1(_06922_),
    .A2(_06926_),
    .A3(_06927_),
    .ZN(_06928_));
 OAI21_X1 _30458_ (.A(_06876_),
    .B1(_06877_),
    .B2(_06920_),
    .ZN(_06929_));
 XNOR2_X2 _30459_ (.A(_06900_),
    .B(_06929_),
    .ZN(_06930_));
 NAND3_X1 _30460_ (.A1(_06919_),
    .A2(_06928_),
    .A3(_06930_),
    .ZN(_06931_));
 INV_X1 _30461_ (.A(_06931_),
    .ZN(_06932_));
 AOI21_X1 _30462_ (.A(_06796_),
    .B1(_19475_),
    .B2(_06801_),
    .ZN(_06933_));
 OAI21_X1 _30463_ (.A(_06826_),
    .B1(_06829_),
    .B2(_06933_),
    .ZN(_06934_));
 AOI21_X1 _30464_ (.A(_06822_),
    .B1(_06825_),
    .B2(_06934_),
    .ZN(_06935_));
 OAI221_X1 _30465_ (.A(_06854_),
    .B1(_06915_),
    .B2(_06916_),
    .C1(_06917_),
    .C2(_06935_),
    .ZN(_06936_));
 AOI21_X1 _30466_ (.A(_19451_),
    .B1(_06936_),
    .B2(_06855_),
    .ZN(_06937_));
 OAI21_X1 _30467_ (.A(_06899_),
    .B1(_06900_),
    .B2(_06937_),
    .ZN(_06938_));
 AOI21_X1 _30468_ (.A(_19447_),
    .B1(_06938_),
    .B2(_06867_),
    .ZN(_06939_));
 OAI21_X1 _30469_ (.A(_06850_),
    .B1(_06851_),
    .B2(_06939_),
    .ZN(_06940_));
 XOR2_X2 _30470_ (.A(_19444_),
    .B(_06940_),
    .Z(_06941_));
 AND4_X1 _30471_ (.A1(_06898_),
    .A2(_06914_),
    .A3(_06932_),
    .A4(_06941_),
    .ZN(_06942_));
 AND2_X1 _30472_ (.A1(_06893_),
    .A2(_06942_),
    .ZN(_06943_));
 XOR2_X1 _30473_ (.A(_06871_),
    .B(_06943_),
    .Z(_14218_));
 INV_X1 _30474_ (.A(_14218_),
    .ZN(_14221_));
 INV_X2 _30475_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.b ),
    .ZN(_06944_));
 CLKBUF_X3 _30476_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.b ),
    .Z(_06945_));
 NOR4_X2 _30477_ (.A1(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_06945_),
    .ZN(_06946_));
 NAND2_X4 _30478_ (.A1(_06944_),
    .A2(_06946_),
    .ZN(_06947_));
 OR4_X1 _30479_ (.A1(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_06948_));
 OAI21_X2 _30480_ (.A(_06947_),
    .B1(_06948_),
    .B2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_06949_));
 NAND4_X2 _30481_ (.A1(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_06945_),
    .ZN(_06950_));
 NOR2_X4 _30482_ (.A1(_06944_),
    .A2(_06950_),
    .ZN(_06951_));
 AND4_X1 _30483_ (.A1(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_06952_));
 AOI21_X4 _30484_ (.A(_06951_),
    .B1(_06952_),
    .B2(\g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_06953_));
 INV_X1 _30485_ (.A(_14220_),
    .ZN(_06954_));
 AOI21_X1 _30486_ (.A(_06949_),
    .B1(_06953_),
    .B2(_06954_),
    .ZN(_00193_));
 INV_X1 _30487_ (.A(_19484_),
    .ZN(_06955_));
 AOI21_X1 _30488_ (.A(_06949_),
    .B1(_06953_),
    .B2(_06955_),
    .ZN(_00194_));
 INV_X1 _30489_ (.A(_14229_),
    .ZN(_06956_));
 AOI21_X1 _30490_ (.A(_06949_),
    .B1(_06953_),
    .B2(_06956_),
    .ZN(_00195_));
 XOR2_X1 _30491_ (.A(_14228_),
    .B(_19493_),
    .Z(_06957_));
 AOI21_X1 _30492_ (.A(_06949_),
    .B1(_06953_),
    .B2(_06957_),
    .ZN(_00196_));
 AOI21_X1 _30493_ (.A(_19488_),
    .B1(_19489_),
    .B2(_19483_),
    .ZN(_06958_));
 INV_X1 _30494_ (.A(_06958_),
    .ZN(_06959_));
 AOI21_X1 _30495_ (.A(_19492_),
    .B1(_06959_),
    .B2(_19493_),
    .ZN(_06960_));
 XNOR2_X1 _30496_ (.A(_06945_),
    .B(_19490_),
    .ZN(_06961_));
 XNOR2_X1 _30497_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_06961_),
    .ZN(_06962_));
 XNOR2_X1 _30498_ (.A(_06960_),
    .B(_06962_),
    .ZN(_06963_));
 AOI21_X1 _30499_ (.A(_06949_),
    .B1(_06953_),
    .B2(_06963_),
    .ZN(_00197_));
 INV_X1 _30500_ (.A(_06949_),
    .ZN(_06964_));
 NAND2_X4 _30501_ (.A1(_06964_),
    .A2(_06953_),
    .ZN(_06965_));
 NAND2_X1 _30502_ (.A1(_19497_),
    .A2(_14218_),
    .ZN(_06966_));
 NAND3_X1 _30503_ (.A1(_06810_),
    .A2(_06847_),
    .A3(_14221_),
    .ZN(_06967_));
 AOI21_X2 _30504_ (.A(_06965_),
    .B1(_06966_),
    .B2(_06967_),
    .ZN(_00192_));
 INV_X1 _30505_ (.A(_19497_),
    .ZN(_06968_));
 XNOR2_X1 _30506_ (.A(_19496_),
    .B(_06921_),
    .ZN(_06969_));
 MUX2_X1 _30507_ (.A(_06968_),
    .B(_06969_),
    .S(_14218_),
    .Z(_06970_));
 NOR2_X1 _30508_ (.A1(_06965_),
    .A2(_06970_),
    .ZN(_00198_));
 XNOR2_X1 _30509_ (.A(_06922_),
    .B(_06927_),
    .ZN(_06971_));
 MUX2_X1 _30510_ (.A(_06969_),
    .B(_06971_),
    .S(_14218_),
    .Z(_06972_));
 NOR2_X1 _30511_ (.A1(_06965_),
    .A2(_06972_),
    .ZN(_00199_));
 NAND3_X1 _30512_ (.A1(_19496_),
    .A2(_06921_),
    .A3(_06927_),
    .ZN(_06973_));
 XNOR2_X1 _30513_ (.A(_06925_),
    .B(_06973_),
    .ZN(_06974_));
 MUX2_X1 _30514_ (.A(_06971_),
    .B(_06974_),
    .S(_14218_),
    .Z(_06975_));
 NOR2_X1 _30515_ (.A1(_06965_),
    .A2(_06975_),
    .ZN(_00200_));
 XNOR2_X1 _30516_ (.A(_06919_),
    .B(_06928_),
    .ZN(_06976_));
 MUX2_X1 _30517_ (.A(_06974_),
    .B(_06976_),
    .S(_14218_),
    .Z(_06977_));
 NOR2_X1 _30518_ (.A1(_06965_),
    .A2(_06977_),
    .ZN(_00201_));
 INV_X1 _30519_ (.A(_06919_),
    .ZN(_06978_));
 NOR3_X1 _30520_ (.A1(_06978_),
    .A2(_06925_),
    .A3(_06973_),
    .ZN(_06979_));
 XNOR2_X1 _30521_ (.A(_06930_),
    .B(_06979_),
    .ZN(_06980_));
 MUX2_X1 _30522_ (.A(_06976_),
    .B(_06980_),
    .S(_14218_),
    .Z(_06981_));
 NOR2_X1 _30523_ (.A1(_06965_),
    .A2(_06981_),
    .ZN(_00202_));
 XOR2_X1 _30524_ (.A(_06898_),
    .B(_06931_),
    .Z(_06982_));
 MUX2_X1 _30525_ (.A(_06980_),
    .B(_06982_),
    .S(_14218_),
    .Z(_06983_));
 NOR2_X1 _30526_ (.A1(_06965_),
    .A2(_06983_),
    .ZN(_00203_));
 INV_X1 _30527_ (.A(_06914_),
    .ZN(_06984_));
 NAND3_X1 _30528_ (.A1(_06898_),
    .A2(_06930_),
    .A3(_06979_),
    .ZN(_06985_));
 XNOR2_X1 _30529_ (.A(_06984_),
    .B(_06985_),
    .ZN(_06986_));
 MUX2_X1 _30530_ (.A(_06982_),
    .B(_06986_),
    .S(_14218_),
    .Z(_06987_));
 NOR2_X1 _30531_ (.A1(_06965_),
    .A2(_06987_),
    .ZN(_00204_));
 AOI21_X1 _30532_ (.A(_06965_),
    .B1(_06986_),
    .B2(_06942_),
    .ZN(_06988_));
 NOR2_X1 _30533_ (.A1(_06943_),
    .A2(_06986_),
    .ZN(_06989_));
 AND3_X1 _30534_ (.A1(_06898_),
    .A2(_06914_),
    .A3(_06932_),
    .ZN(_06990_));
 NOR2_X1 _30535_ (.A1(_06990_),
    .A2(_06941_),
    .ZN(_06991_));
 INV_X1 _30536_ (.A(_06893_),
    .ZN(_06992_));
 AOI21_X1 _30537_ (.A(_06991_),
    .B1(_06942_),
    .B2(_06992_),
    .ZN(_06993_));
 MUX2_X1 _30538_ (.A(_06989_),
    .B(_06993_),
    .S(_06871_),
    .Z(_06994_));
 AND2_X1 _30539_ (.A1(_06988_),
    .A2(_06994_),
    .ZN(_00205_));
 NOR2_X1 _30540_ (.A1(_06984_),
    .A2(_06985_),
    .ZN(_06995_));
 NAND4_X1 _30541_ (.A1(_06871_),
    .A2(_06992_),
    .A3(_06941_),
    .A4(_06995_),
    .ZN(_06996_));
 OAI21_X1 _30542_ (.A(_06941_),
    .B1(_06995_),
    .B2(_06990_),
    .ZN(_06997_));
 NOR2_X1 _30543_ (.A1(_06871_),
    .A2(_06995_),
    .ZN(_06998_));
 AOI22_X2 _30544_ (.A1(_06871_),
    .A2(_06997_),
    .B1(_06998_),
    .B2(_06990_),
    .ZN(_06999_));
 XNOR2_X1 _30545_ (.A(_06990_),
    .B(_06941_),
    .ZN(_07000_));
 OAI221_X1 _30546_ (.A(_06996_),
    .B1(_06999_),
    .B2(_06992_),
    .C1(_06871_),
    .C2(_07000_),
    .ZN(_07001_));
 AND3_X1 _30547_ (.A1(_06964_),
    .A2(_06953_),
    .A3(_07001_),
    .ZN(_00206_));
 CLKBUF_X2 _30548_ (.A(_19523_),
    .Z(_07002_));
 INV_X1 _30549_ (.A(_07002_),
    .ZN(_07003_));
 INV_X1 _30550_ (.A(_19524_),
    .ZN(_07004_));
 CLKBUF_X2 _30551_ (.A(_19527_),
    .Z(_07005_));
 INV_X1 _30552_ (.A(_19528_),
    .ZN(_07006_));
 BUF_X1 _30553_ (.A(_19530_),
    .Z(_07007_));
 INV_X1 _30554_ (.A(_19532_),
    .ZN(_07008_));
 AOI21_X1 _30555_ (.A(_19534_),
    .B1(_19535_),
    .B2(_19536_),
    .ZN(_07009_));
 INV_X1 _30556_ (.A(_19533_),
    .ZN(_07010_));
 OAI21_X1 _30557_ (.A(_07008_),
    .B1(_07009_),
    .B2(_07010_),
    .ZN(_07011_));
 BUF_X1 _30558_ (.A(_19531_),
    .Z(_07012_));
 AOI21_X1 _30559_ (.A(_07007_),
    .B1(_07011_),
    .B2(_07012_),
    .ZN(_07013_));
 INV_X1 _30560_ (.A(_19529_),
    .ZN(_07014_));
 OAI21_X1 _30561_ (.A(_07006_),
    .B1(_07013_),
    .B2(_07014_),
    .ZN(_07015_));
 AOI21_X1 _30562_ (.A(_19526_),
    .B1(_07005_),
    .B2(_07015_),
    .ZN(_07016_));
 CLKBUF_X2 _30563_ (.A(_19525_),
    .Z(_07017_));
 INV_X1 _30564_ (.A(_07017_),
    .ZN(_07018_));
 OAI21_X1 _30565_ (.A(_07004_),
    .B1(_07016_),
    .B2(_07018_),
    .ZN(_07019_));
 XNOR2_X1 _30566_ (.A(_07003_),
    .B(_07019_),
    .ZN(_07020_));
 CLKBUF_X2 _30567_ (.A(_19521_),
    .Z(_07021_));
 INV_X1 _30568_ (.A(_07021_),
    .ZN(_07022_));
 AOI21_X1 _30569_ (.A(_19522_),
    .B1(_07002_),
    .B2(_19524_),
    .ZN(_07023_));
 NAND2_X1 _30570_ (.A1(_07002_),
    .A2(_07017_),
    .ZN(_07024_));
 AOI21_X2 _30571_ (.A(_19526_),
    .B1(_07005_),
    .B2(_19528_),
    .ZN(_07025_));
 OAI21_X1 _30572_ (.A(_07023_),
    .B1(_07024_),
    .B2(_07025_),
    .ZN(_07026_));
 INV_X1 _30573_ (.A(_07026_),
    .ZN(_07027_));
 OAI21_X1 _30574_ (.A(_07008_),
    .B1(_07010_),
    .B2(_14233_),
    .ZN(_07028_));
 AOI21_X1 _30575_ (.A(_07007_),
    .B1(_07028_),
    .B2(_07012_),
    .ZN(_07029_));
 NAND2_X1 _30576_ (.A1(_07005_),
    .A2(_19529_),
    .ZN(_07030_));
 OR2_X1 _30577_ (.A1(_07029_),
    .A2(_07030_),
    .ZN(_07031_));
 OAI21_X1 _30578_ (.A(_07027_),
    .B1(_07031_),
    .B2(_07024_),
    .ZN(_07032_));
 XNOR2_X1 _30579_ (.A(_07022_),
    .B(_07032_),
    .ZN(_07033_));
 XNOR2_X1 _30580_ (.A(_14233_),
    .B(_19533_),
    .ZN(_07034_));
 NOR4_X1 _30581_ (.A1(_14234_),
    .A2(\g_row[0].g_col[1].mult.adder.a[0] ),
    .A3(_19537_),
    .A4(_07034_),
    .ZN(_07035_));
 XNOR2_X1 _30582_ (.A(_07014_),
    .B(_07029_),
    .ZN(_07036_));
 XNOR2_X1 _30583_ (.A(_07012_),
    .B(_07011_),
    .ZN(_07037_));
 AND2_X1 _30584_ (.A1(_07025_),
    .A2(_07031_),
    .ZN(_07038_));
 XNOR2_X1 _30585_ (.A(_07018_),
    .B(_07038_),
    .ZN(_07039_));
 NAND4_X1 _30586_ (.A1(_07035_),
    .A2(_07036_),
    .A3(_07037_),
    .A4(_07039_),
    .ZN(_07040_));
 XNOR2_X1 _30587_ (.A(_07005_),
    .B(_07015_),
    .ZN(_07041_));
 BUF_X2 _30588_ (.A(_19517_),
    .Z(_07042_));
 BUF_X2 _30589_ (.A(_19519_),
    .Z(_07043_));
 INV_X1 _30590_ (.A(_19520_),
    .ZN(_07044_));
 OAI21_X1 _30591_ (.A(_07044_),
    .B1(_07023_),
    .B2(_07022_),
    .ZN(_07045_));
 AOI21_X1 _30592_ (.A(_19518_),
    .B1(_07043_),
    .B2(_07045_),
    .ZN(_07046_));
 NAND4_X2 _30593_ (.A1(_07043_),
    .A2(_07021_),
    .A3(_07002_),
    .A4(_07017_),
    .ZN(_07047_));
 OAI21_X2 _30594_ (.A(_07046_),
    .B1(_07047_),
    .B2(_07038_),
    .ZN(_07048_));
 XNOR2_X2 _30595_ (.A(_07042_),
    .B(_07048_),
    .ZN(_07049_));
 NAND2_X1 _30596_ (.A1(_07041_),
    .A2(_07049_),
    .ZN(_07050_));
 NOR4_X2 _30597_ (.A1(_07020_),
    .A2(_07033_),
    .A3(_07040_),
    .A4(_07050_),
    .ZN(_07051_));
 AOI21_X1 _30598_ (.A(_19522_),
    .B1(_07002_),
    .B2(_07019_),
    .ZN(_07052_));
 OAI21_X1 _30599_ (.A(_07044_),
    .B1(_07052_),
    .B2(_07022_),
    .ZN(_07053_));
 XNOR2_X2 _30600_ (.A(_07043_),
    .B(_07053_),
    .ZN(_07054_));
 NOR2_X1 _30601_ (.A1(_07051_),
    .A2(_07054_),
    .ZN(_19551_));
 INV_X1 _30602_ (.A(_19498_),
    .ZN(_07055_));
 INV_X1 _30603_ (.A(_19499_),
    .ZN(_07056_));
 INV_X1 _30604_ (.A(_19502_),
    .ZN(_07057_));
 INV_X2 _30605_ (.A(_19503_),
    .ZN(_07058_));
 BUF_X1 _30606_ (.A(_19504_),
    .Z(_07059_));
 BUF_X1 _30607_ (.A(_19506_),
    .Z(_07060_));
 CLKBUF_X2 _30608_ (.A(_19507_),
    .Z(_07061_));
 INV_X1 _30609_ (.A(_19508_),
    .ZN(_07062_));
 BUF_X2 _30610_ (.A(_19511_),
    .Z(_07063_));
 AOI21_X1 _30611_ (.A(_19510_),
    .B1(_07063_),
    .B2(_19512_),
    .ZN(_07064_));
 BUF_X2 _30612_ (.A(_19509_),
    .Z(_07065_));
 INV_X1 _30613_ (.A(_07065_),
    .ZN(_07066_));
 OAI21_X1 _30614_ (.A(_07062_),
    .B1(_07064_),
    .B2(_07066_),
    .ZN(_07067_));
 AOI21_X1 _30615_ (.A(_07060_),
    .B1(_07061_),
    .B2(_07067_),
    .ZN(_07068_));
 BUF_X2 _30616_ (.A(_19515_),
    .Z(_07069_));
 AOI21_X1 _30617_ (.A(_19514_),
    .B1(_07069_),
    .B2(_19516_),
    .ZN(_07070_));
 INV_X1 _30618_ (.A(_19518_),
    .ZN(_07071_));
 INV_X1 _30619_ (.A(_07043_),
    .ZN(_07072_));
 AOI21_X1 _30620_ (.A(_19520_),
    .B1(_07026_),
    .B2(_07021_),
    .ZN(_07073_));
 OAI21_X1 _30621_ (.A(_07071_),
    .B1(_07072_),
    .B2(_07073_),
    .ZN(_07074_));
 NAND3_X1 _30622_ (.A1(_07069_),
    .A2(_07042_),
    .A3(_07074_),
    .ZN(_07075_));
 AND2_X1 _30623_ (.A1(_07070_),
    .A2(_07075_),
    .ZN(_07076_));
 BUF_X2 _30624_ (.A(_19513_),
    .Z(_07077_));
 NAND4_X1 _30625_ (.A1(_07061_),
    .A2(_07065_),
    .A3(_07063_),
    .A4(_07077_),
    .ZN(_07078_));
 OAI21_X1 _30626_ (.A(_07068_),
    .B1(_07076_),
    .B2(_07078_),
    .ZN(_07079_));
 BUF_X2 _30627_ (.A(_19505_),
    .Z(_07080_));
 AOI21_X1 _30628_ (.A(_07059_),
    .B1(_07079_),
    .B2(_07080_),
    .ZN(_07081_));
 OAI21_X1 _30629_ (.A(_07057_),
    .B1(_07058_),
    .B2(_07081_),
    .ZN(_07082_));
 AOI21_X1 _30630_ (.A(_19500_),
    .B1(_19501_),
    .B2(_07082_),
    .ZN(_07083_));
 OAI21_X2 _30631_ (.A(_07055_),
    .B1(_07056_),
    .B2(_07083_),
    .ZN(_07084_));
 INV_X1 _30632_ (.A(_19510_),
    .ZN(_07085_));
 INV_X1 _30633_ (.A(_07063_),
    .ZN(_07086_));
 AOI21_X1 _30634_ (.A(_19512_),
    .B1(_07077_),
    .B2(_19514_),
    .ZN(_07087_));
 OAI21_X1 _30635_ (.A(_07085_),
    .B1(_07086_),
    .B2(_07087_),
    .ZN(_07088_));
 AOI21_X1 _30636_ (.A(_19508_),
    .B1(_07088_),
    .B2(_07065_),
    .ZN(_07089_));
 AND2_X1 _30637_ (.A1(_07077_),
    .A2(_07069_),
    .ZN(_07090_));
 NAND3_X1 _30638_ (.A1(_07065_),
    .A2(_07063_),
    .A3(_07090_),
    .ZN(_07091_));
 INV_X1 _30639_ (.A(_19522_),
    .ZN(_07092_));
 INV_X1 _30640_ (.A(_19526_),
    .ZN(_07093_));
 INV_X1 _30641_ (.A(_07005_),
    .ZN(_07094_));
 AOI21_X1 _30642_ (.A(_19528_),
    .B1(_07007_),
    .B2(_19529_),
    .ZN(_07095_));
 OAI21_X1 _30643_ (.A(_07093_),
    .B1(_07094_),
    .B2(_07095_),
    .ZN(_07096_));
 AOI21_X1 _30644_ (.A(_19524_),
    .B1(_07096_),
    .B2(_07017_),
    .ZN(_07097_));
 OAI21_X1 _30645_ (.A(_07092_),
    .B1(_07003_),
    .B2(_07097_),
    .ZN(_07098_));
 AOI21_X1 _30646_ (.A(_19520_),
    .B1(_07098_),
    .B2(_07021_),
    .ZN(_07099_));
 OAI21_X1 _30647_ (.A(_07071_),
    .B1(_07072_),
    .B2(_07099_),
    .ZN(_07100_));
 AOI21_X1 _30648_ (.A(_19516_),
    .B1(_07100_),
    .B2(_07042_),
    .ZN(_07101_));
 OAI21_X1 _30649_ (.A(_07089_),
    .B1(_07091_),
    .B2(_07101_),
    .ZN(_07102_));
 AOI21_X1 _30650_ (.A(_07060_),
    .B1(_07061_),
    .B2(_07102_),
    .ZN(_07103_));
 INV_X1 _30651_ (.A(_07103_),
    .ZN(_07104_));
 AOI21_X1 _30652_ (.A(_07059_),
    .B1(_07104_),
    .B2(_07080_),
    .ZN(_07105_));
 OAI21_X1 _30653_ (.A(_07057_),
    .B1(_07058_),
    .B2(_07105_),
    .ZN(_07106_));
 AOI21_X2 _30654_ (.A(_19500_),
    .B1(_19501_),
    .B2(_07106_),
    .ZN(_07107_));
 XNOR2_X2 _30655_ (.A(_19499_),
    .B(_07107_),
    .ZN(_07108_));
 OR3_X1 _30656_ (.A1(_07060_),
    .A2(_07058_),
    .A3(_07059_),
    .ZN(_07109_));
 NAND2_X1 _30657_ (.A1(_07077_),
    .A2(_07069_),
    .ZN(_07110_));
 INV_X1 _30658_ (.A(_07007_),
    .ZN(_07111_));
 AOI21_X1 _30659_ (.A(_19532_),
    .B1(_19534_),
    .B2(_19533_),
    .ZN(_07112_));
 INV_X1 _30660_ (.A(_07012_),
    .ZN(_07113_));
 OAI21_X1 _30661_ (.A(_07111_),
    .B1(_07112_),
    .B2(_07113_),
    .ZN(_07114_));
 AOI21_X1 _30662_ (.A(_19528_),
    .B1(_07114_),
    .B2(_19529_),
    .ZN(_07115_));
 OAI21_X1 _30663_ (.A(_07093_),
    .B1(_07094_),
    .B2(_07115_),
    .ZN(_07116_));
 AOI21_X1 _30664_ (.A(_19524_),
    .B1(_07116_),
    .B2(_07017_),
    .ZN(_07117_));
 OAI21_X1 _30665_ (.A(_07092_),
    .B1(_07003_),
    .B2(_07117_),
    .ZN(_07118_));
 AOI21_X1 _30666_ (.A(_19520_),
    .B1(_07118_),
    .B2(_07021_),
    .ZN(_07119_));
 OAI21_X1 _30667_ (.A(_07071_),
    .B1(_07072_),
    .B2(_07119_),
    .ZN(_07120_));
 AOI21_X1 _30668_ (.A(_19516_),
    .B1(_07120_),
    .B2(_07042_),
    .ZN(_07121_));
 OAI21_X1 _30669_ (.A(_07087_),
    .B1(_07110_),
    .B2(_07121_),
    .ZN(_07122_));
 AOI21_X1 _30670_ (.A(_19510_),
    .B1(_07063_),
    .B2(_07122_),
    .ZN(_07123_));
 OAI21_X1 _30671_ (.A(_07062_),
    .B1(_07123_),
    .B2(_07066_),
    .ZN(_07124_));
 AOI21_X2 _30672_ (.A(_07109_),
    .B1(_07124_),
    .B2(_07061_),
    .ZN(_07125_));
 AND4_X1 _30673_ (.A1(_07058_),
    .A2(_07080_),
    .A3(_07061_),
    .A4(_07124_),
    .ZN(_07126_));
 NAND2_X1 _30674_ (.A1(_07058_),
    .A2(_07059_),
    .ZN(_07127_));
 OR3_X1 _30675_ (.A1(_07058_),
    .A2(_07080_),
    .A3(_07059_),
    .ZN(_07128_));
 NAND3_X1 _30676_ (.A1(_07060_),
    .A2(_07058_),
    .A3(_07080_),
    .ZN(_07129_));
 NAND3_X2 _30677_ (.A1(_07127_),
    .A2(_07128_),
    .A3(_07129_),
    .ZN(_07130_));
 NOR3_X4 _30678_ (.A1(_07125_),
    .A2(_07126_),
    .A3(_07130_),
    .ZN(_07131_));
 NAND2_X1 _30679_ (.A1(_07069_),
    .A2(_07042_),
    .ZN(_07132_));
 OR3_X1 _30680_ (.A1(_07031_),
    .A2(_07047_),
    .A3(_07132_),
    .ZN(_07133_));
 AND2_X1 _30681_ (.A1(_07076_),
    .A2(_07133_),
    .ZN(_07134_));
 OAI21_X1 _30682_ (.A(_07068_),
    .B1(_07078_),
    .B2(_07134_),
    .ZN(_07135_));
 XNOR2_X2 _30683_ (.A(_07080_),
    .B(_07135_),
    .ZN(_07136_));
 INV_X1 _30684_ (.A(_19516_),
    .ZN(_07137_));
 AOI21_X1 _30685_ (.A(_19518_),
    .B1(_07043_),
    .B2(_07053_),
    .ZN(_07138_));
 INV_X1 _30686_ (.A(_07042_),
    .ZN(_07139_));
 OAI21_X1 _30687_ (.A(_07137_),
    .B1(_07138_),
    .B2(_07139_),
    .ZN(_07140_));
 AOI221_X2 _30688_ (.A(_19512_),
    .B1(_07090_),
    .B2(_07140_),
    .C1(_07077_),
    .C2(_19514_),
    .ZN(_07141_));
 XNOR2_X2 _30689_ (.A(_07063_),
    .B(_07141_),
    .ZN(_07142_));
 XNOR2_X1 _30690_ (.A(_07069_),
    .B(_07140_),
    .ZN(_07143_));
 NOR3_X1 _30691_ (.A1(_07049_),
    .A2(_07054_),
    .A3(_07143_),
    .ZN(_07144_));
 XNOR2_X2 _30692_ (.A(_07077_),
    .B(_07134_),
    .ZN(_07145_));
 AND3_X1 _30693_ (.A1(_07142_),
    .A2(_07144_),
    .A3(_07145_),
    .ZN(_07146_));
 NAND2_X1 _30694_ (.A1(_07063_),
    .A2(_07077_),
    .ZN(_07147_));
 OAI21_X1 _30695_ (.A(_07064_),
    .B1(_07070_),
    .B2(_07147_),
    .ZN(_07148_));
 NOR2_X1 _30696_ (.A1(_07132_),
    .A2(_07147_),
    .ZN(_07149_));
 AOI21_X2 _30697_ (.A(_07148_),
    .B1(_07149_),
    .B2(_07048_),
    .ZN(_07150_));
 XNOR2_X2 _30698_ (.A(_07065_),
    .B(_07150_),
    .ZN(_07151_));
 INV_X1 _30699_ (.A(_07061_),
    .ZN(_07152_));
 NAND4_X1 _30700_ (.A1(_07065_),
    .A2(_07063_),
    .A3(_07090_),
    .A4(_07140_),
    .ZN(_07153_));
 NAND2_X1 _30701_ (.A1(_07089_),
    .A2(_07153_),
    .ZN(_07154_));
 XNOR2_X1 _30702_ (.A(_07152_),
    .B(_07154_),
    .ZN(_07155_));
 NAND3_X1 _30703_ (.A1(_07146_),
    .A2(_07151_),
    .A3(_07155_),
    .ZN(_07156_));
 OR3_X1 _30704_ (.A1(_07131_),
    .A2(_07136_),
    .A3(_07156_),
    .ZN(_07157_));
 INV_X1 _30705_ (.A(_07059_),
    .ZN(_07158_));
 NOR3_X1 _30706_ (.A1(_07072_),
    .A2(_07022_),
    .A3(_07024_),
    .ZN(_07159_));
 AOI21_X1 _30707_ (.A(_07007_),
    .B1(_19532_),
    .B2(_07012_),
    .ZN(_07160_));
 OAI21_X1 _30708_ (.A(_07025_),
    .B1(_07030_),
    .B2(_07160_),
    .ZN(_07161_));
 AOI221_X2 _30709_ (.A(_19518_),
    .B1(_07043_),
    .B2(_07045_),
    .C1(_07159_),
    .C2(_07161_),
    .ZN(_07162_));
 NOR3_X1 _30710_ (.A1(_07132_),
    .A2(_07147_),
    .A3(_07162_),
    .ZN(_07163_));
 OAI21_X1 _30711_ (.A(_07065_),
    .B1(_07148_),
    .B2(_07163_),
    .ZN(_07164_));
 AOI21_X1 _30712_ (.A(_07152_),
    .B1(_07062_),
    .B2(_07164_),
    .ZN(_07165_));
 OAI21_X1 _30713_ (.A(_07080_),
    .B1(_07165_),
    .B2(_07060_),
    .ZN(_07166_));
 AOI21_X1 _30714_ (.A(_07058_),
    .B1(_07158_),
    .B2(_07166_),
    .ZN(_07167_));
 NOR2_X1 _30715_ (.A1(_19502_),
    .A2(_07167_),
    .ZN(_07168_));
 XNOR2_X2 _30716_ (.A(_19501_),
    .B(_07168_),
    .ZN(_07169_));
 INV_X1 _30717_ (.A(_07169_),
    .ZN(_07170_));
 NOR2_X1 _30718_ (.A1(_07157_),
    .A2(_07170_),
    .ZN(_07171_));
 NAND2_X1 _30719_ (.A1(_07108_),
    .A2(_07171_),
    .ZN(_07172_));
 XNOR2_X1 _30720_ (.A(_07084_),
    .B(_07172_),
    .ZN(_14237_));
 INV_X1 _30721_ (.A(_14237_),
    .ZN(_14240_));
 INV_X2 _30722_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.b ),
    .ZN(_07173_));
 BUF_X4 _30723_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.b ),
    .Z(_07174_));
 NOR4_X2 _30724_ (.A1(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07174_),
    .ZN(_07175_));
 NAND2_X4 _30725_ (.A1(_07173_),
    .A2(_07175_),
    .ZN(_07176_));
 OR4_X1 _30726_ (.A1(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07177_));
 OAI21_X2 _30727_ (.A(_07176_),
    .B1(_07177_),
    .B2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07178_));
 NAND4_X2 _30728_ (.A1(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07174_),
    .ZN(_07179_));
 NOR2_X4 _30729_ (.A1(_07173_),
    .A2(_07179_),
    .ZN(_07180_));
 AND4_X1 _30730_ (.A1(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07181_));
 AOI21_X4 _30731_ (.A(_07180_),
    .B1(_07181_),
    .B2(\g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07182_));
 INV_X1 _30732_ (.A(_14239_),
    .ZN(_07183_));
 AOI21_X1 _30733_ (.A(_07178_),
    .B1(_07182_),
    .B2(_07183_),
    .ZN(_00209_));
 INV_X1 _30734_ (.A(_19541_),
    .ZN(_07184_));
 AOI21_X1 _30735_ (.A(_07178_),
    .B1(_07182_),
    .B2(_07184_),
    .ZN(_00210_));
 INV_X1 _30736_ (.A(_14248_),
    .ZN(_07185_));
 AOI21_X1 _30737_ (.A(_07178_),
    .B1(_07182_),
    .B2(_07185_),
    .ZN(_00211_));
 XOR2_X1 _30738_ (.A(_14247_),
    .B(_19550_),
    .Z(_07186_));
 AOI21_X1 _30739_ (.A(_07178_),
    .B1(_07182_),
    .B2(_07186_),
    .ZN(_00212_));
 AOI21_X1 _30740_ (.A(_19545_),
    .B1(_19546_),
    .B2(_19540_),
    .ZN(_07187_));
 INV_X1 _30741_ (.A(_07187_),
    .ZN(_07188_));
 AOI21_X1 _30742_ (.A(_19549_),
    .B1(_07188_),
    .B2(_19550_),
    .ZN(_07189_));
 XNOR2_X1 _30743_ (.A(_07174_),
    .B(_19547_),
    .ZN(_07190_));
 XNOR2_X1 _30744_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_07190_),
    .ZN(_07191_));
 XNOR2_X1 _30745_ (.A(_07189_),
    .B(_07191_),
    .ZN(_07192_));
 AOI21_X1 _30746_ (.A(_07178_),
    .B1(_07182_),
    .B2(_07192_),
    .ZN(_00213_));
 INV_X1 _30747_ (.A(_07178_),
    .ZN(_07193_));
 NAND2_X4 _30748_ (.A1(_07193_),
    .A2(_07182_),
    .ZN(_07194_));
 INV_X1 _30749_ (.A(_07194_),
    .ZN(_07195_));
 NAND2_X1 _30750_ (.A1(_07051_),
    .A2(_07195_),
    .ZN(_07196_));
 NOR2_X1 _30751_ (.A1(_07054_),
    .A2(_07196_),
    .ZN(_07197_));
 AND2_X1 _30752_ (.A1(_19554_),
    .A2(_07195_),
    .ZN(_07198_));
 MUX2_X1 _30753_ (.A(_07197_),
    .B(_07198_),
    .S(_14237_),
    .Z(_00208_));
 XOR2_X1 _30754_ (.A(_19553_),
    .B(_07143_),
    .Z(_07199_));
 NOR2_X1 _30755_ (.A1(_07194_),
    .A2(_07199_),
    .ZN(_07200_));
 MUX2_X1 _30756_ (.A(_07198_),
    .B(_07200_),
    .S(_14237_),
    .Z(_00214_));
 XNOR2_X1 _30757_ (.A(_07144_),
    .B(_07145_),
    .ZN(_07201_));
 NOR2_X1 _30758_ (.A1(_07194_),
    .A2(_07201_),
    .ZN(_07202_));
 MUX2_X1 _30759_ (.A(_07200_),
    .B(_07202_),
    .S(_14237_),
    .Z(_00215_));
 NAND2_X1 _30760_ (.A1(_19553_),
    .A2(_07145_),
    .ZN(_07203_));
 NOR2_X1 _30761_ (.A1(_07143_),
    .A2(_07203_),
    .ZN(_07204_));
 XNOR2_X1 _30762_ (.A(_07142_),
    .B(_07204_),
    .ZN(_07205_));
 NOR2_X1 _30763_ (.A1(_07194_),
    .A2(_07205_),
    .ZN(_07206_));
 MUX2_X1 _30764_ (.A(_07202_),
    .B(_07206_),
    .S(_14237_),
    .Z(_00216_));
 XNOR2_X1 _30765_ (.A(_07146_),
    .B(_07151_),
    .ZN(_07207_));
 NOR2_X1 _30766_ (.A1(_07194_),
    .A2(_07207_),
    .ZN(_07208_));
 MUX2_X1 _30767_ (.A(_07206_),
    .B(_07208_),
    .S(_14237_),
    .Z(_00217_));
 INV_X1 _30768_ (.A(_07155_),
    .ZN(_07209_));
 NAND3_X1 _30769_ (.A1(_07142_),
    .A2(_07151_),
    .A3(_07204_),
    .ZN(_07210_));
 XNOR2_X1 _30770_ (.A(_07209_),
    .B(_07210_),
    .ZN(_07211_));
 NOR2_X1 _30771_ (.A1(_07194_),
    .A2(_07211_),
    .ZN(_07212_));
 MUX2_X1 _30772_ (.A(_07208_),
    .B(_07212_),
    .S(_14237_),
    .Z(_00218_));
 XNOR2_X1 _30773_ (.A(_07136_),
    .B(_07156_),
    .ZN(_07213_));
 NOR2_X1 _30774_ (.A1(_07194_),
    .A2(_07213_),
    .ZN(_07214_));
 MUX2_X1 _30775_ (.A(_07212_),
    .B(_07214_),
    .S(_14237_),
    .Z(_00219_));
 OR3_X2 _30776_ (.A1(_07136_),
    .A2(_07209_),
    .A3(_07210_),
    .ZN(_07215_));
 XNOR2_X2 _30777_ (.A(_07131_),
    .B(_07215_),
    .ZN(_07216_));
 NOR2_X1 _30778_ (.A1(_07194_),
    .A2(_07216_),
    .ZN(_07217_));
 MUX2_X1 _30779_ (.A(_07214_),
    .B(_07217_),
    .S(_14237_),
    .Z(_00220_));
 AOI21_X1 _30780_ (.A(_07194_),
    .B1(_07216_),
    .B2(_07171_),
    .ZN(_07218_));
 AOI21_X1 _30781_ (.A(_07216_),
    .B1(_07171_),
    .B2(_07108_),
    .ZN(_07219_));
 INV_X1 _30782_ (.A(_07157_),
    .ZN(_07220_));
 NOR2_X1 _30783_ (.A1(_07220_),
    .A2(_07169_),
    .ZN(_07221_));
 INV_X1 _30784_ (.A(_07108_),
    .ZN(_07222_));
 AOI21_X1 _30785_ (.A(_07221_),
    .B1(_07171_),
    .B2(_07222_),
    .ZN(_07223_));
 MUX2_X1 _30786_ (.A(_07219_),
    .B(_07223_),
    .S(_07084_),
    .Z(_07224_));
 AND2_X1 _30787_ (.A1(_07218_),
    .A2(_07224_),
    .ZN(_00221_));
 OAI21_X1 _30788_ (.A(_07108_),
    .B1(_07215_),
    .B2(_07131_),
    .ZN(_07225_));
 AOI21_X1 _30789_ (.A(_07221_),
    .B1(_07225_),
    .B2(_07171_),
    .ZN(_07226_));
 NOR2_X1 _30790_ (.A1(_07131_),
    .A2(_07215_),
    .ZN(_07227_));
 OAI21_X1 _30791_ (.A(_07169_),
    .B1(_07227_),
    .B2(_07220_),
    .ZN(_07228_));
 NOR3_X1 _30792_ (.A1(_07131_),
    .A2(_07170_),
    .A3(_07215_),
    .ZN(_07229_));
 MUX2_X1 _30793_ (.A(_07228_),
    .B(_07229_),
    .S(_07222_),
    .Z(_07230_));
 MUX2_X1 _30794_ (.A(_07226_),
    .B(_07230_),
    .S(_07084_),
    .Z(_07231_));
 AND2_X1 _30795_ (.A1(_07195_),
    .A2(_07231_),
    .ZN(_00222_));
 BUF_X2 _30796_ (.A(_19578_),
    .Z(_07232_));
 AOI21_X2 _30797_ (.A(_19577_),
    .B1(_07232_),
    .B2(_19579_),
    .ZN(_07233_));
 CLKBUF_X2 _30798_ (.A(_19580_),
    .Z(_07234_));
 NAND2_X2 _30799_ (.A1(_07232_),
    .A2(_07234_),
    .ZN(_07235_));
 CLKBUF_X2 _30800_ (.A(_19583_),
    .Z(_07236_));
 AOI21_X1 _30801_ (.A(_19581_),
    .B1(_19582_),
    .B2(_07236_),
    .ZN(_07237_));
 OAI21_X1 _30802_ (.A(_07233_),
    .B1(_07235_),
    .B2(_07237_),
    .ZN(_07238_));
 INV_X1 _30803_ (.A(_19582_),
    .ZN(_07239_));
 NOR2_X1 _30804_ (.A1(_07239_),
    .A2(_07235_),
    .ZN(_07240_));
 BUF_X2 _30805_ (.A(_19584_),
    .Z(_07241_));
 INV_X1 _30806_ (.A(_19585_),
    .ZN(_07242_));
 CLKBUF_X2 _30807_ (.A(_19587_),
    .Z(_07243_));
 INV_X1 _30808_ (.A(_19589_),
    .ZN(_07244_));
 AOI21_X1 _30809_ (.A(_19591_),
    .B1(_19592_),
    .B2(_19593_),
    .ZN(_07245_));
 INV_X1 _30810_ (.A(_19590_),
    .ZN(_07246_));
 OAI21_X1 _30811_ (.A(_07244_),
    .B1(_07245_),
    .B2(_07246_),
    .ZN(_07247_));
 AOI21_X1 _30812_ (.A(_07243_),
    .B1(_07247_),
    .B2(_19588_),
    .ZN(_07248_));
 BUF_X1 _30813_ (.A(_19586_),
    .Z(_07249_));
 INV_X1 _30814_ (.A(_07249_),
    .ZN(_07250_));
 OAI21_X1 _30815_ (.A(_07242_),
    .B1(_07248_),
    .B2(_07250_),
    .ZN(_07251_));
 AND2_X1 _30816_ (.A1(_07241_),
    .A2(_07251_),
    .ZN(_07252_));
 AOI21_X2 _30817_ (.A(_07238_),
    .B1(_07240_),
    .B2(_07252_),
    .ZN(_07253_));
 XNOR2_X1 _30818_ (.A(_19576_),
    .B(_07253_),
    .ZN(_07254_));
 INV_X1 _30819_ (.A(_19581_),
    .ZN(_07255_));
 OAI21_X1 _30820_ (.A(_19582_),
    .B1(_07252_),
    .B2(_07236_),
    .ZN(_07256_));
 NAND2_X1 _30821_ (.A1(_07255_),
    .A2(_07256_),
    .ZN(_07257_));
 XOR2_X1 _30822_ (.A(_07234_),
    .B(_07257_),
    .Z(_07258_));
 BUF_X2 _30823_ (.A(_19574_),
    .Z(_07259_));
 INV_X1 _30824_ (.A(_19575_),
    .ZN(_07260_));
 INV_X1 _30825_ (.A(_19576_),
    .ZN(_07261_));
 AOI21_X1 _30826_ (.A(_19579_),
    .B1(_07234_),
    .B2(_19581_),
    .ZN(_07262_));
 INV_X1 _30827_ (.A(_07262_),
    .ZN(_07263_));
 AOI21_X1 _30828_ (.A(_19577_),
    .B1(_07263_),
    .B2(_07232_),
    .ZN(_07264_));
 OAI21_X1 _30829_ (.A(_07260_),
    .B1(_07261_),
    .B2(_07264_),
    .ZN(_07265_));
 NOR3_X2 _30830_ (.A1(_07261_),
    .A2(_07239_),
    .A3(_07235_),
    .ZN(_07266_));
 AOI21_X2 _30831_ (.A(_07236_),
    .B1(_07241_),
    .B2(_19585_),
    .ZN(_07267_));
 OAI21_X1 _30832_ (.A(_07244_),
    .B1(_07246_),
    .B2(_14252_),
    .ZN(_07268_));
 AOI21_X2 _30833_ (.A(_07243_),
    .B1(_07268_),
    .B2(_19588_),
    .ZN(_07269_));
 NAND2_X1 _30834_ (.A1(_07241_),
    .A2(_07249_),
    .ZN(_07270_));
 OAI21_X1 _30835_ (.A(_07267_),
    .B1(_07269_),
    .B2(_07270_),
    .ZN(_07271_));
 AOI21_X2 _30836_ (.A(_07265_),
    .B1(_07266_),
    .B2(_07271_),
    .ZN(_07272_));
 XNOR2_X2 _30837_ (.A(_07259_),
    .B(_07272_),
    .ZN(_19608_));
 XOR2_X1 _30838_ (.A(_07241_),
    .B(_07251_),
    .Z(_07273_));
 NAND2_X1 _30839_ (.A1(_07250_),
    .A2(_07242_),
    .ZN(_07274_));
 AOI21_X1 _30840_ (.A(_07236_),
    .B1(_07241_),
    .B2(_07274_),
    .ZN(_07275_));
 XNOR2_X1 _30841_ (.A(_07239_),
    .B(_07275_),
    .ZN(_07276_));
 XNOR2_X1 _30842_ (.A(_14252_),
    .B(_19590_),
    .ZN(_07277_));
 NOR4_X1 _30843_ (.A1(_14253_),
    .A2(\g_row[0].g_col[2].mult.adder.a[0] ),
    .A3(_19594_),
    .A4(_07277_),
    .ZN(_07278_));
 NAND2_X1 _30844_ (.A1(_07239_),
    .A2(_07255_),
    .ZN(_07279_));
 AOI21_X1 _30845_ (.A(_19579_),
    .B1(_07234_),
    .B2(_07279_),
    .ZN(_07280_));
 XOR2_X1 _30846_ (.A(_07232_),
    .B(_07280_),
    .Z(_07281_));
 XNOR2_X1 _30847_ (.A(_07249_),
    .B(_07269_),
    .ZN(_07282_));
 INV_X1 _30848_ (.A(_19588_),
    .ZN(_07283_));
 XNOR2_X1 _30849_ (.A(_07283_),
    .B(_07247_),
    .ZN(_07284_));
 NOR2_X1 _30850_ (.A1(_07282_),
    .A2(_07284_),
    .ZN(_07285_));
 NAND4_X1 _30851_ (.A1(_07276_),
    .A2(_07278_),
    .A3(_07281_),
    .A4(_07285_),
    .ZN(_07286_));
 OR4_X1 _30852_ (.A1(_07258_),
    .A2(_19608_),
    .A3(_07273_),
    .A4(_07286_),
    .ZN(_07287_));
 AND2_X1 _30853_ (.A1(_07254_),
    .A2(_07287_),
    .ZN(_19609_));
 INV_X1 _30854_ (.A(_19555_),
    .ZN(_07288_));
 INV_X1 _30855_ (.A(_19556_),
    .ZN(_07289_));
 INV_X1 _30856_ (.A(_19559_),
    .ZN(_07290_));
 INV_X1 _30857_ (.A(_19560_),
    .ZN(_07291_));
 INV_X1 _30858_ (.A(_19565_),
    .ZN(_07292_));
 BUF_X2 _30859_ (.A(_19568_),
    .Z(_07293_));
 AOI21_X2 _30860_ (.A(_19567_),
    .B1(_07293_),
    .B2(_19569_),
    .ZN(_07294_));
 CLKBUF_X2 _30861_ (.A(_19566_),
    .Z(_07295_));
 INV_X1 _30862_ (.A(_07295_),
    .ZN(_07296_));
 OAI21_X1 _30863_ (.A(_07292_),
    .B1(_07294_),
    .B2(_07296_),
    .ZN(_07297_));
 AOI21_X1 _30864_ (.A(_19563_),
    .B1(_19564_),
    .B2(_07297_),
    .ZN(_07298_));
 BUF_X2 _30865_ (.A(_19572_),
    .Z(_07299_));
 BUF_X2 _30866_ (.A(_19573_),
    .Z(_07300_));
 AND2_X1 _30867_ (.A1(_07299_),
    .A2(_07259_),
    .ZN(_07301_));
 NAND2_X1 _30868_ (.A1(_07234_),
    .A2(_19582_),
    .ZN(_07302_));
 OAI21_X1 _30869_ (.A(_07262_),
    .B1(_07267_),
    .B2(_07302_),
    .ZN(_07303_));
 AOI21_X1 _30870_ (.A(_19577_),
    .B1(_07303_),
    .B2(_07232_),
    .ZN(_07304_));
 OAI21_X1 _30871_ (.A(_07260_),
    .B1(_07261_),
    .B2(_07304_),
    .ZN(_07305_));
 AOI221_X2 _30872_ (.A(_19571_),
    .B1(_07299_),
    .B2(_07300_),
    .C1(_07301_),
    .C2(_07305_),
    .ZN(_07306_));
 BUF_X2 _30873_ (.A(_19570_),
    .Z(_07307_));
 NAND4_X1 _30874_ (.A1(_19564_),
    .A2(_07295_),
    .A3(_07293_),
    .A4(_07307_),
    .ZN(_07308_));
 OAI21_X1 _30875_ (.A(_07298_),
    .B1(_07306_),
    .B2(_07308_),
    .ZN(_07309_));
 BUF_X2 _30876_ (.A(_19562_),
    .Z(_07310_));
 AOI21_X1 _30877_ (.A(_19561_),
    .B1(_07309_),
    .B2(_07310_),
    .ZN(_07311_));
 OAI21_X1 _30878_ (.A(_07290_),
    .B1(_07291_),
    .B2(_07311_),
    .ZN(_07312_));
 AOI21_X2 _30879_ (.A(_19557_),
    .B1(_19558_),
    .B2(_07312_),
    .ZN(_07313_));
 OAI21_X4 _30880_ (.A(_07288_),
    .B1(_07289_),
    .B2(_07313_),
    .ZN(_07314_));
 INV_X1 _30881_ (.A(_19563_),
    .ZN(_07315_));
 INV_X1 _30882_ (.A(_19564_),
    .ZN(_07316_));
 AOI21_X2 _30883_ (.A(_19571_),
    .B1(_07299_),
    .B2(_07300_),
    .ZN(_07317_));
 NAND2_X1 _30884_ (.A1(_07293_),
    .A2(_07307_),
    .ZN(_07318_));
 NAND3_X1 _30885_ (.A1(_07293_),
    .A2(_07307_),
    .A3(_07301_),
    .ZN(_07319_));
 AOI21_X1 _30886_ (.A(_07243_),
    .B1(_19589_),
    .B2(_19588_),
    .ZN(_07320_));
 OAI21_X1 _30887_ (.A(_07267_),
    .B1(_07270_),
    .B2(_07320_),
    .ZN(_07321_));
 AOI21_X1 _30888_ (.A(_07265_),
    .B1(_07266_),
    .B2(_07321_),
    .ZN(_07322_));
 OAI221_X1 _30889_ (.A(_07294_),
    .B1(_07317_),
    .B2(_07318_),
    .C1(_07319_),
    .C2(_07322_),
    .ZN(_07323_));
 AOI21_X1 _30890_ (.A(_19565_),
    .B1(_07323_),
    .B2(_07295_),
    .ZN(_07324_));
 OAI21_X1 _30891_ (.A(_07315_),
    .B1(_07316_),
    .B2(_07324_),
    .ZN(_07325_));
 AOI21_X1 _30892_ (.A(_19561_),
    .B1(_07325_),
    .B2(_07310_),
    .ZN(_07326_));
 OAI21_X1 _30893_ (.A(_07290_),
    .B1(_07291_),
    .B2(_07326_),
    .ZN(_07327_));
 XNOR2_X2 _30894_ (.A(_19558_),
    .B(_07327_),
    .ZN(_07328_));
 INV_X1 _30895_ (.A(_19567_),
    .ZN(_07329_));
 INV_X1 _30896_ (.A(_07293_),
    .ZN(_07330_));
 AOI21_X1 _30897_ (.A(_19569_),
    .B1(_07307_),
    .B2(_19571_),
    .ZN(_07331_));
 OAI21_X1 _30898_ (.A(_07329_),
    .B1(_07330_),
    .B2(_07331_),
    .ZN(_07332_));
 AOI21_X1 _30899_ (.A(_19565_),
    .B1(_07332_),
    .B2(_07295_),
    .ZN(_07333_));
 NAND4_X1 _30900_ (.A1(_07295_),
    .A2(_07293_),
    .A3(_07307_),
    .A4(_07299_),
    .ZN(_07334_));
 NAND2_X1 _30901_ (.A1(_07259_),
    .A2(_19576_),
    .ZN(_07335_));
 NOR2_X1 _30902_ (.A1(_07235_),
    .A2(_07335_),
    .ZN(_07336_));
 AOI21_X1 _30903_ (.A(_19585_),
    .B1(_07243_),
    .B2(_07249_),
    .ZN(_07337_));
 INV_X1 _30904_ (.A(_07337_),
    .ZN(_07338_));
 AOI21_X1 _30905_ (.A(_07236_),
    .B1(_07241_),
    .B2(_07338_),
    .ZN(_07339_));
 OAI21_X1 _30906_ (.A(_07255_),
    .B1(_07339_),
    .B2(_07239_),
    .ZN(_07340_));
 OAI21_X2 _30907_ (.A(_07260_),
    .B1(_07261_),
    .B2(_07233_),
    .ZN(_07341_));
 AOI221_X2 _30908_ (.A(_07300_),
    .B1(_07336_),
    .B2(_07340_),
    .C1(_07341_),
    .C2(_07259_),
    .ZN(_07342_));
 OAI21_X1 _30909_ (.A(_07333_),
    .B1(_07334_),
    .B2(_07342_),
    .ZN(_07343_));
 AOI21_X1 _30910_ (.A(_19563_),
    .B1(_19564_),
    .B2(_07343_),
    .ZN(_07344_));
 INV_X1 _30911_ (.A(_07344_),
    .ZN(_07345_));
 AOI21_X1 _30912_ (.A(_19561_),
    .B1(_07345_),
    .B2(_07310_),
    .ZN(_07346_));
 OAI21_X1 _30913_ (.A(_07290_),
    .B1(_07291_),
    .B2(_07346_),
    .ZN(_07347_));
 AOI21_X2 _30914_ (.A(_19557_),
    .B1(_19558_),
    .B2(_07347_),
    .ZN(_07348_));
 XNOR2_X2 _30915_ (.A(_19556_),
    .B(_07348_),
    .ZN(_07349_));
 INV_X1 _30916_ (.A(_07349_),
    .ZN(_07350_));
 NOR2_X1 _30917_ (.A1(_07269_),
    .A2(_07270_),
    .ZN(_07351_));
 NAND3_X1 _30918_ (.A1(_07266_),
    .A2(_07351_),
    .A3(_07301_),
    .ZN(_07352_));
 NAND2_X1 _30919_ (.A1(_07306_),
    .A2(_07352_),
    .ZN(_07353_));
 INV_X1 _30920_ (.A(_07353_),
    .ZN(_07354_));
 OAI21_X1 _30921_ (.A(_07298_),
    .B1(_07308_),
    .B2(_07354_),
    .ZN(_07355_));
 XOR2_X2 _30922_ (.A(_07310_),
    .B(_07355_),
    .Z(_07356_));
 NAND2_X1 _30923_ (.A1(_07307_),
    .A2(_07299_),
    .ZN(_07357_));
 AOI21_X1 _30924_ (.A(_07300_),
    .B1(_07259_),
    .B2(_19575_),
    .ZN(_07358_));
 OAI21_X1 _30925_ (.A(_07331_),
    .B1(_07357_),
    .B2(_07358_),
    .ZN(_07359_));
 NOR2_X1 _30926_ (.A1(_07357_),
    .A2(_07335_),
    .ZN(_07360_));
 NAND2_X1 _30927_ (.A1(_07241_),
    .A2(_07240_),
    .ZN(_07361_));
 INV_X1 _30928_ (.A(_07243_),
    .ZN(_07362_));
 AOI21_X1 _30929_ (.A(_19589_),
    .B1(_19591_),
    .B2(_19590_),
    .ZN(_07363_));
 OAI21_X1 _30930_ (.A(_07362_),
    .B1(_07363_),
    .B2(_07283_),
    .ZN(_07364_));
 AOI21_X1 _30931_ (.A(_19585_),
    .B1(_07364_),
    .B2(_07249_),
    .ZN(_07365_));
 OAI221_X1 _30932_ (.A(_07233_),
    .B1(_07235_),
    .B2(_07237_),
    .C1(_07361_),
    .C2(_07365_),
    .ZN(_07366_));
 AOI21_X1 _30933_ (.A(_07359_),
    .B1(_07360_),
    .B2(_07366_),
    .ZN(_07367_));
 OAI21_X1 _30934_ (.A(_07329_),
    .B1(_07330_),
    .B2(_07367_),
    .ZN(_07368_));
 AOI21_X1 _30935_ (.A(_19565_),
    .B1(_07368_),
    .B2(_07295_),
    .ZN(_07369_));
 OAI21_X1 _30936_ (.A(_07315_),
    .B1(_07316_),
    .B2(_07369_),
    .ZN(_07370_));
 AOI21_X2 _30937_ (.A(_19561_),
    .B1(_07370_),
    .B2(_07310_),
    .ZN(_07371_));
 XNOR2_X2 _30938_ (.A(_19560_),
    .B(_07371_),
    .ZN(_07372_));
 OAI221_X2 _30939_ (.A(_07294_),
    .B1(_07317_),
    .B2(_07318_),
    .C1(_07319_),
    .C2(_07272_),
    .ZN(_07373_));
 XNOR2_X2 _30940_ (.A(_07296_),
    .B(_07373_),
    .ZN(_07374_));
 AOI221_X1 _30941_ (.A(_07300_),
    .B1(_07257_),
    .B2(_07336_),
    .C1(_07341_),
    .C2(_07259_),
    .ZN(_07375_));
 XNOR2_X2 _30942_ (.A(_07299_),
    .B(_07375_),
    .ZN(_07376_));
 AND3_X1 _30943_ (.A1(_07254_),
    .A2(_19608_),
    .A3(_07376_),
    .ZN(_07377_));
 NOR3_X1 _30944_ (.A1(_07253_),
    .A2(_07357_),
    .A3(_07335_),
    .ZN(_07378_));
 NOR2_X1 _30945_ (.A1(_07359_),
    .A2(_07378_),
    .ZN(_07379_));
 XNOR2_X2 _30946_ (.A(_07330_),
    .B(_07379_),
    .ZN(_07380_));
 INV_X1 _30947_ (.A(_07380_),
    .ZN(_07381_));
 XOR2_X2 _30948_ (.A(_07307_),
    .B(_07353_),
    .Z(_07382_));
 AND3_X1 _30949_ (.A1(_07377_),
    .A2(_07381_),
    .A3(_07382_),
    .ZN(_07383_));
 OAI21_X1 _30950_ (.A(_07333_),
    .B1(_07334_),
    .B2(_07375_),
    .ZN(_07384_));
 XNOR2_X2 _30951_ (.A(_07316_),
    .B(_07384_),
    .ZN(_07385_));
 NAND3_X1 _30952_ (.A1(_07374_),
    .A2(_07383_),
    .A3(_07385_),
    .ZN(_07386_));
 INV_X1 _30953_ (.A(_07386_),
    .ZN(_07387_));
 NAND3_X1 _30954_ (.A1(_07356_),
    .A2(_07372_),
    .A3(_07387_),
    .ZN(_07388_));
 NOR3_X1 _30955_ (.A1(_07328_),
    .A2(_07350_),
    .A3(_07388_),
    .ZN(_07389_));
 XOR2_X2 _30956_ (.A(_07314_),
    .B(_07389_),
    .Z(_07390_));
 BUF_X1 _30957_ (.A(_07390_),
    .Z(_14256_));
 INV_X1 _30958_ (.A(_14256_),
    .ZN(_14261_));
 INV_X2 _30959_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.b ),
    .ZN(_07391_));
 CLKBUF_X3 _30960_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.b ),
    .Z(_07392_));
 NOR4_X2 _30961_ (.A1(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07392_),
    .ZN(_07393_));
 NAND2_X4 _30962_ (.A1(_07391_),
    .A2(_07393_),
    .ZN(_07394_));
 OR4_X2 _30963_ (.A1(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07395_));
 OAI21_X4 _30964_ (.A(_07394_),
    .B1(_07395_),
    .B2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07396_));
 NAND4_X2 _30965_ (.A1(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07392_),
    .ZN(_07397_));
 NOR2_X4 _30966_ (.A1(_07391_),
    .A2(_07397_),
    .ZN(_07398_));
 AND4_X1 _30967_ (.A1(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07399_));
 AOI21_X4 _30968_ (.A(_07398_),
    .B1(_07399_),
    .B2(\g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07400_));
 INV_X1 _30969_ (.A(_14258_),
    .ZN(_07401_));
 AOI21_X1 _30970_ (.A(_07396_),
    .B1(_07400_),
    .B2(_07401_),
    .ZN(_00225_));
 INV_X1 _30971_ (.A(_19598_),
    .ZN(_07402_));
 AOI21_X1 _30972_ (.A(_07396_),
    .B1(_07400_),
    .B2(_07402_),
    .ZN(_00226_));
 INV_X1 _30973_ (.A(_14267_),
    .ZN(_07403_));
 AOI21_X1 _30974_ (.A(_07396_),
    .B1(_07400_),
    .B2(_07403_),
    .ZN(_00227_));
 XOR2_X1 _30975_ (.A(_14266_),
    .B(_19607_),
    .Z(_07404_));
 AOI21_X1 _30976_ (.A(_07396_),
    .B1(_07400_),
    .B2(_07404_),
    .ZN(_00228_));
 AOI21_X1 _30977_ (.A(_19602_),
    .B1(_19603_),
    .B2(_19597_),
    .ZN(_07405_));
 INV_X1 _30978_ (.A(_07405_),
    .ZN(_07406_));
 AOI21_X1 _30979_ (.A(_19606_),
    .B1(_07406_),
    .B2(_19607_),
    .ZN(_07407_));
 XNOR2_X1 _30980_ (.A(_07392_),
    .B(_19604_),
    .ZN(_07408_));
 XNOR2_X1 _30981_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_07408_),
    .ZN(_07409_));
 XNOR2_X1 _30982_ (.A(_07407_),
    .B(_07409_),
    .ZN(_07410_));
 AOI21_X1 _30983_ (.A(_07396_),
    .B1(_07400_),
    .B2(_07410_),
    .ZN(_00229_));
 INV_X1 _30984_ (.A(_07396_),
    .ZN(_07411_));
 NAND2_X4 _30985_ (.A1(_07411_),
    .A2(_07400_),
    .ZN(_07412_));
 INV_X1 _30986_ (.A(_07287_),
    .ZN(_07413_));
 NAND2_X1 _30987_ (.A1(_07254_),
    .A2(_07413_),
    .ZN(_07414_));
 INV_X1 _30988_ (.A(_19611_),
    .ZN(_07415_));
 MUX2_X1 _30989_ (.A(_07414_),
    .B(_07415_),
    .S(_14256_),
    .Z(_07416_));
 NOR2_X1 _30990_ (.A1(_07412_),
    .A2(_07416_),
    .ZN(_00224_));
 XNOR2_X1 _30991_ (.A(_19610_),
    .B(_07376_),
    .ZN(_07417_));
 MUX2_X1 _30992_ (.A(_07415_),
    .B(_07417_),
    .S(_14256_),
    .Z(_07418_));
 NOR2_X2 _30993_ (.A1(_07412_),
    .A2(_07418_),
    .ZN(_00230_));
 XNOR2_X1 _30994_ (.A(_07377_),
    .B(_07382_),
    .ZN(_07419_));
 MUX2_X1 _30995_ (.A(_07417_),
    .B(_07419_),
    .S(_14256_),
    .Z(_07420_));
 NOR2_X1 _30996_ (.A1(_07412_),
    .A2(_07420_),
    .ZN(_00231_));
 NAND3_X1 _30997_ (.A1(_19610_),
    .A2(_07376_),
    .A3(_07382_),
    .ZN(_07421_));
 XNOR2_X1 _30998_ (.A(_07380_),
    .B(_07421_),
    .ZN(_07422_));
 MUX2_X1 _30999_ (.A(_07419_),
    .B(_07422_),
    .S(_14256_),
    .Z(_07423_));
 NOR2_X1 _31000_ (.A1(_07412_),
    .A2(_07423_),
    .ZN(_00232_));
 XNOR2_X1 _31001_ (.A(_07374_),
    .B(_07383_),
    .ZN(_07424_));
 MUX2_X1 _31002_ (.A(_07422_),
    .B(_07424_),
    .S(_14256_),
    .Z(_07425_));
 NOR2_X1 _31003_ (.A1(_07412_),
    .A2(_07425_),
    .ZN(_00233_));
 INV_X1 _31004_ (.A(_07374_),
    .ZN(_07426_));
 NOR3_X1 _31005_ (.A1(_07426_),
    .A2(_07380_),
    .A3(_07421_),
    .ZN(_07427_));
 XNOR2_X1 _31006_ (.A(_07385_),
    .B(_07427_),
    .ZN(_07428_));
 MUX2_X1 _31007_ (.A(_07424_),
    .B(_07428_),
    .S(_14256_),
    .Z(_07429_));
 NOR2_X1 _31008_ (.A1(_07412_),
    .A2(_07429_),
    .ZN(_00234_));
 XOR2_X1 _31009_ (.A(_07356_),
    .B(_07386_),
    .Z(_07430_));
 MUX2_X1 _31010_ (.A(_07428_),
    .B(_07430_),
    .S(_14256_),
    .Z(_07431_));
 NOR2_X1 _31011_ (.A1(_07412_),
    .A2(_07431_),
    .ZN(_00235_));
 NAND3_X1 _31012_ (.A1(_07356_),
    .A2(_07385_),
    .A3(_07427_),
    .ZN(_07432_));
 XOR2_X1 _31013_ (.A(_07372_),
    .B(_07432_),
    .Z(_07433_));
 MUX2_X1 _31014_ (.A(_07430_),
    .B(_07433_),
    .S(_14256_),
    .Z(_07434_));
 NOR2_X1 _31015_ (.A1(_07412_),
    .A2(_07434_),
    .ZN(_00236_));
 XNOR2_X1 _31016_ (.A(_07328_),
    .B(_07388_),
    .ZN(_07435_));
 MUX2_X1 _31017_ (.A(_07433_),
    .B(_07435_),
    .S(_07390_),
    .Z(_07436_));
 NOR2_X1 _31018_ (.A1(_07412_),
    .A2(_07436_),
    .ZN(_00237_));
 NAND4_X2 _31019_ (.A1(_07356_),
    .A2(_07372_),
    .A3(_07385_),
    .A4(_07427_),
    .ZN(_07437_));
 NAND4_X1 _31020_ (.A1(_07314_),
    .A2(_07349_),
    .A3(_07388_),
    .A4(_07437_),
    .ZN(_07438_));
 AOI21_X1 _31021_ (.A(_07388_),
    .B1(_07437_),
    .B2(_07349_),
    .ZN(_07439_));
 NOR2_X1 _31022_ (.A1(_07314_),
    .A2(_07439_),
    .ZN(_07440_));
 NOR2_X1 _31023_ (.A1(_07349_),
    .A2(_07437_),
    .ZN(_07441_));
 AOI21_X1 _31024_ (.A(_07440_),
    .B1(_07441_),
    .B2(_07314_),
    .ZN(_07442_));
 NAND2_X1 _31025_ (.A1(_07314_),
    .A2(_07349_),
    .ZN(_07443_));
 OAI21_X1 _31026_ (.A(_07443_),
    .B1(_07388_),
    .B2(_07314_),
    .ZN(_07444_));
 INV_X1 _31027_ (.A(_07444_),
    .ZN(_07445_));
 MUX2_X1 _31028_ (.A(_07442_),
    .B(_07445_),
    .S(_07328_),
    .Z(_07446_));
 AOI21_X2 _31029_ (.A(_07412_),
    .B1(_07438_),
    .B2(_07446_),
    .ZN(_00238_));
 CLKBUF_X2 _31030_ (.A(_19637_),
    .Z(_07447_));
 INV_X1 _31031_ (.A(_07447_),
    .ZN(_07448_));
 INV_X1 _31032_ (.A(_19638_),
    .ZN(_07449_));
 CLKBUF_X2 _31033_ (.A(_19641_),
    .Z(_07450_));
 INV_X1 _31034_ (.A(_19642_),
    .ZN(_07451_));
 BUF_X1 _31035_ (.A(_19644_),
    .Z(_07452_));
 INV_X1 _31036_ (.A(_19646_),
    .ZN(_07453_));
 AOI21_X1 _31037_ (.A(_19648_),
    .B1(_19649_),
    .B2(_19650_),
    .ZN(_07454_));
 INV_X1 _31038_ (.A(_19647_),
    .ZN(_07455_));
 OAI21_X1 _31039_ (.A(_07453_),
    .B1(_07454_),
    .B2(_07455_),
    .ZN(_07456_));
 BUF_X1 _31040_ (.A(_19645_),
    .Z(_07457_));
 AOI21_X1 _31041_ (.A(_07452_),
    .B1(_07456_),
    .B2(_07457_),
    .ZN(_07458_));
 INV_X1 _31042_ (.A(_19643_),
    .ZN(_07459_));
 OAI21_X1 _31043_ (.A(_07451_),
    .B1(_07458_),
    .B2(_07459_),
    .ZN(_07460_));
 AOI21_X1 _31044_ (.A(_19640_),
    .B1(_07450_),
    .B2(_07460_),
    .ZN(_07461_));
 CLKBUF_X2 _31045_ (.A(_19639_),
    .Z(_07462_));
 INV_X1 _31046_ (.A(_07462_),
    .ZN(_07463_));
 OAI21_X1 _31047_ (.A(_07449_),
    .B1(_07461_),
    .B2(_07463_),
    .ZN(_07464_));
 XNOR2_X1 _31048_ (.A(_07448_),
    .B(_07464_),
    .ZN(_07465_));
 CLKBUF_X2 _31049_ (.A(_19635_),
    .Z(_07466_));
 INV_X1 _31050_ (.A(_07466_),
    .ZN(_07467_));
 AOI21_X1 _31051_ (.A(_19636_),
    .B1(_07447_),
    .B2(_19638_),
    .ZN(_07468_));
 NAND2_X1 _31052_ (.A1(_07447_),
    .A2(_07462_),
    .ZN(_07469_));
 AOI21_X2 _31053_ (.A(_19640_),
    .B1(_07450_),
    .B2(_19642_),
    .ZN(_07470_));
 OAI21_X1 _31054_ (.A(_07468_),
    .B1(_07469_),
    .B2(_07470_),
    .ZN(_07471_));
 INV_X1 _31055_ (.A(_07471_),
    .ZN(_07472_));
 OAI21_X1 _31056_ (.A(_07453_),
    .B1(_07455_),
    .B2(_14271_),
    .ZN(_07473_));
 AOI21_X1 _31057_ (.A(_07452_),
    .B1(_07473_),
    .B2(_07457_),
    .ZN(_07474_));
 NAND2_X1 _31058_ (.A1(_07450_),
    .A2(_19643_),
    .ZN(_07475_));
 OR2_X1 _31059_ (.A1(_07474_),
    .A2(_07475_),
    .ZN(_07476_));
 OAI21_X1 _31060_ (.A(_07472_),
    .B1(_07476_),
    .B2(_07469_),
    .ZN(_07477_));
 XNOR2_X1 _31061_ (.A(_07467_),
    .B(_07477_),
    .ZN(_07478_));
 XNOR2_X1 _31062_ (.A(_14271_),
    .B(_19647_),
    .ZN(_07479_));
 NOR4_X1 _31063_ (.A1(_14272_),
    .A2(\g_row[0].g_col[3].mult.adder.a[0] ),
    .A3(_19651_),
    .A4(_07479_),
    .ZN(_07480_));
 XNOR2_X1 _31064_ (.A(_07459_),
    .B(_07474_),
    .ZN(_07481_));
 XNOR2_X1 _31065_ (.A(_07457_),
    .B(_07456_),
    .ZN(_07482_));
 AND2_X1 _31066_ (.A1(_07470_),
    .A2(_07476_),
    .ZN(_07483_));
 XNOR2_X1 _31067_ (.A(_07463_),
    .B(_07483_),
    .ZN(_07484_));
 NAND4_X1 _31068_ (.A1(_07480_),
    .A2(_07481_),
    .A3(_07482_),
    .A4(_07484_),
    .ZN(_07485_));
 XNOR2_X1 _31069_ (.A(_07450_),
    .B(_07460_),
    .ZN(_07486_));
 BUF_X2 _31070_ (.A(_19631_),
    .Z(_07487_));
 BUF_X2 _31071_ (.A(_19633_),
    .Z(_07488_));
 INV_X1 _31072_ (.A(_19634_),
    .ZN(_07489_));
 OAI21_X1 _31073_ (.A(_07489_),
    .B1(_07468_),
    .B2(_07467_),
    .ZN(_07490_));
 AOI21_X1 _31074_ (.A(_19632_),
    .B1(_07488_),
    .B2(_07490_),
    .ZN(_07491_));
 NAND4_X2 _31075_ (.A1(_07488_),
    .A2(_07466_),
    .A3(_07447_),
    .A4(_07462_),
    .ZN(_07492_));
 OAI21_X2 _31076_ (.A(_07491_),
    .B1(_07492_),
    .B2(_07483_),
    .ZN(_07493_));
 XNOR2_X2 _31077_ (.A(_07487_),
    .B(_07493_),
    .ZN(_07494_));
 NAND2_X1 _31078_ (.A1(_07486_),
    .A2(_07494_),
    .ZN(_07495_));
 NOR4_X2 _31079_ (.A1(_07465_),
    .A2(_07478_),
    .A3(_07485_),
    .A4(_07495_),
    .ZN(_07496_));
 AOI21_X1 _31080_ (.A(_19636_),
    .B1(_07447_),
    .B2(_07464_),
    .ZN(_07497_));
 OAI21_X1 _31081_ (.A(_07489_),
    .B1(_07497_),
    .B2(_07467_),
    .ZN(_07498_));
 XNOR2_X2 _31082_ (.A(_07488_),
    .B(_07498_),
    .ZN(_07499_));
 NOR2_X1 _31083_ (.A1(_07496_),
    .A2(_07499_),
    .ZN(_19666_));
 INV_X1 _31084_ (.A(_19612_),
    .ZN(_07500_));
 INV_X1 _31085_ (.A(_19613_),
    .ZN(_07501_));
 INV_X1 _31086_ (.A(_19616_),
    .ZN(_07502_));
 INV_X2 _31087_ (.A(_19617_),
    .ZN(_07503_));
 BUF_X1 _31088_ (.A(_19618_),
    .Z(_07504_));
 BUF_X1 _31089_ (.A(_19620_),
    .Z(_07505_));
 CLKBUF_X2 _31090_ (.A(_19621_),
    .Z(_07506_));
 INV_X1 _31091_ (.A(_19622_),
    .ZN(_07507_));
 BUF_X2 _31092_ (.A(_19625_),
    .Z(_07508_));
 AOI21_X1 _31093_ (.A(_19624_),
    .B1(_07508_),
    .B2(_19626_),
    .ZN(_07509_));
 BUF_X2 _31094_ (.A(_19623_),
    .Z(_07510_));
 INV_X1 _31095_ (.A(_07510_),
    .ZN(_07511_));
 OAI21_X1 _31096_ (.A(_07507_),
    .B1(_07509_),
    .B2(_07511_),
    .ZN(_07512_));
 AOI21_X1 _31097_ (.A(_07505_),
    .B1(_07506_),
    .B2(_07512_),
    .ZN(_07513_));
 BUF_X2 _31098_ (.A(_19629_),
    .Z(_07514_));
 AOI21_X1 _31099_ (.A(_19628_),
    .B1(_07514_),
    .B2(_19630_),
    .ZN(_07515_));
 INV_X1 _31100_ (.A(_19632_),
    .ZN(_07516_));
 INV_X1 _31101_ (.A(_07488_),
    .ZN(_07517_));
 AOI21_X1 _31102_ (.A(_19634_),
    .B1(_07471_),
    .B2(_07466_),
    .ZN(_07518_));
 OAI21_X1 _31103_ (.A(_07516_),
    .B1(_07517_),
    .B2(_07518_),
    .ZN(_07519_));
 NAND3_X1 _31104_ (.A1(_07514_),
    .A2(_07487_),
    .A3(_07519_),
    .ZN(_07520_));
 AND2_X1 _31105_ (.A1(_07515_),
    .A2(_07520_),
    .ZN(_07521_));
 BUF_X2 _31106_ (.A(_19627_),
    .Z(_07522_));
 NAND4_X1 _31107_ (.A1(_07506_),
    .A2(_07510_),
    .A3(_07508_),
    .A4(_07522_),
    .ZN(_07523_));
 OAI21_X1 _31108_ (.A(_07513_),
    .B1(_07521_),
    .B2(_07523_),
    .ZN(_07524_));
 CLKBUF_X2 _31109_ (.A(_19619_),
    .Z(_07525_));
 AOI21_X1 _31110_ (.A(_07504_),
    .B1(_07524_),
    .B2(_07525_),
    .ZN(_07526_));
 OAI21_X1 _31111_ (.A(_07502_),
    .B1(_07503_),
    .B2(_07526_),
    .ZN(_07527_));
 AOI21_X1 _31112_ (.A(_19614_),
    .B1(_19615_),
    .B2(_07527_),
    .ZN(_07528_));
 OAI21_X2 _31113_ (.A(_07500_),
    .B1(_07501_),
    .B2(_07528_),
    .ZN(_07529_));
 INV_X1 _31114_ (.A(_19624_),
    .ZN(_07530_));
 INV_X1 _31115_ (.A(_07508_),
    .ZN(_07531_));
 AOI21_X1 _31116_ (.A(_19626_),
    .B1(_07522_),
    .B2(_19628_),
    .ZN(_07532_));
 OAI21_X1 _31117_ (.A(_07530_),
    .B1(_07531_),
    .B2(_07532_),
    .ZN(_07533_));
 AOI21_X1 _31118_ (.A(_19622_),
    .B1(_07533_),
    .B2(_07510_),
    .ZN(_07534_));
 AND2_X1 _31119_ (.A1(_07522_),
    .A2(_07514_),
    .ZN(_07535_));
 NAND3_X1 _31120_ (.A1(_07510_),
    .A2(_07508_),
    .A3(_07535_),
    .ZN(_07536_));
 INV_X1 _31121_ (.A(_19636_),
    .ZN(_07537_));
 INV_X1 _31122_ (.A(_19640_),
    .ZN(_07538_));
 INV_X1 _31123_ (.A(_07450_),
    .ZN(_07539_));
 AOI21_X1 _31124_ (.A(_19642_),
    .B1(_07452_),
    .B2(_19643_),
    .ZN(_07540_));
 OAI21_X1 _31125_ (.A(_07538_),
    .B1(_07539_),
    .B2(_07540_),
    .ZN(_07541_));
 AOI21_X1 _31126_ (.A(_19638_),
    .B1(_07541_),
    .B2(_07462_),
    .ZN(_07542_));
 OAI21_X1 _31127_ (.A(_07537_),
    .B1(_07448_),
    .B2(_07542_),
    .ZN(_07543_));
 AOI21_X1 _31128_ (.A(_19634_),
    .B1(_07543_),
    .B2(_07466_),
    .ZN(_07544_));
 OAI21_X1 _31129_ (.A(_07516_),
    .B1(_07517_),
    .B2(_07544_),
    .ZN(_07545_));
 AOI21_X1 _31130_ (.A(_19630_),
    .B1(_07545_),
    .B2(_07487_),
    .ZN(_07546_));
 OAI21_X1 _31131_ (.A(_07534_),
    .B1(_07536_),
    .B2(_07546_),
    .ZN(_07547_));
 AOI21_X1 _31132_ (.A(_07505_),
    .B1(_07506_),
    .B2(_07547_),
    .ZN(_07548_));
 INV_X1 _31133_ (.A(_07548_),
    .ZN(_07549_));
 AOI21_X1 _31134_ (.A(_07504_),
    .B1(_07549_),
    .B2(_07525_),
    .ZN(_07550_));
 OAI21_X1 _31135_ (.A(_07502_),
    .B1(_07503_),
    .B2(_07550_),
    .ZN(_07551_));
 AOI21_X2 _31136_ (.A(_19614_),
    .B1(_19615_),
    .B2(_07551_),
    .ZN(_07552_));
 XNOR2_X2 _31137_ (.A(_19613_),
    .B(_07552_),
    .ZN(_07553_));
 OR3_X1 _31138_ (.A1(_07505_),
    .A2(_07503_),
    .A3(_07504_),
    .ZN(_07554_));
 NAND2_X1 _31139_ (.A1(_07522_),
    .A2(_07514_),
    .ZN(_07555_));
 INV_X1 _31140_ (.A(_07452_),
    .ZN(_07556_));
 AOI21_X1 _31141_ (.A(_19646_),
    .B1(_19648_),
    .B2(_19647_),
    .ZN(_07557_));
 INV_X1 _31142_ (.A(_07457_),
    .ZN(_07558_));
 OAI21_X1 _31143_ (.A(_07556_),
    .B1(_07557_),
    .B2(_07558_),
    .ZN(_07559_));
 AOI21_X1 _31144_ (.A(_19642_),
    .B1(_07559_),
    .B2(_19643_),
    .ZN(_07560_));
 OAI21_X1 _31145_ (.A(_07538_),
    .B1(_07539_),
    .B2(_07560_),
    .ZN(_07561_));
 AOI21_X1 _31146_ (.A(_19638_),
    .B1(_07561_),
    .B2(_07462_),
    .ZN(_07562_));
 OAI21_X1 _31147_ (.A(_07537_),
    .B1(_07448_),
    .B2(_07562_),
    .ZN(_07563_));
 AOI21_X1 _31148_ (.A(_19634_),
    .B1(_07563_),
    .B2(_07466_),
    .ZN(_07564_));
 OAI21_X1 _31149_ (.A(_07516_),
    .B1(_07517_),
    .B2(_07564_),
    .ZN(_07565_));
 AOI21_X1 _31150_ (.A(_19630_),
    .B1(_07565_),
    .B2(_07487_),
    .ZN(_07566_));
 OAI21_X1 _31151_ (.A(_07532_),
    .B1(_07555_),
    .B2(_07566_),
    .ZN(_07567_));
 AOI21_X1 _31152_ (.A(_19624_),
    .B1(_07508_),
    .B2(_07567_),
    .ZN(_07568_));
 OAI21_X1 _31153_ (.A(_07507_),
    .B1(_07568_),
    .B2(_07511_),
    .ZN(_07569_));
 AOI21_X2 _31154_ (.A(_07554_),
    .B1(_07569_),
    .B2(_07506_),
    .ZN(_07570_));
 AND4_X1 _31155_ (.A1(_07503_),
    .A2(_07525_),
    .A3(_07506_),
    .A4(_07569_),
    .ZN(_07571_));
 NAND2_X1 _31156_ (.A1(_07503_),
    .A2(_07504_),
    .ZN(_07572_));
 OR3_X1 _31157_ (.A1(_07503_),
    .A2(_07525_),
    .A3(_07504_),
    .ZN(_07573_));
 NAND3_X1 _31158_ (.A1(_07505_),
    .A2(_07503_),
    .A3(_07525_),
    .ZN(_07574_));
 NAND3_X2 _31159_ (.A1(_07572_),
    .A2(_07573_),
    .A3(_07574_),
    .ZN(_07575_));
 NOR3_X4 _31160_ (.A1(_07570_),
    .A2(_07571_),
    .A3(_07575_),
    .ZN(_07576_));
 NAND2_X1 _31161_ (.A1(_07514_),
    .A2(_07487_),
    .ZN(_07577_));
 OR3_X1 _31162_ (.A1(_07476_),
    .A2(_07492_),
    .A3(_07577_),
    .ZN(_07578_));
 AND2_X1 _31163_ (.A1(_07521_),
    .A2(_07578_),
    .ZN(_07579_));
 OAI21_X1 _31164_ (.A(_07513_),
    .B1(_07523_),
    .B2(_07579_),
    .ZN(_07580_));
 XNOR2_X1 _31165_ (.A(_07525_),
    .B(_07580_),
    .ZN(_07581_));
 INV_X1 _31166_ (.A(_19630_),
    .ZN(_07582_));
 AOI21_X1 _31167_ (.A(_19632_),
    .B1(_07488_),
    .B2(_07498_),
    .ZN(_07583_));
 INV_X1 _31168_ (.A(_07487_),
    .ZN(_07584_));
 OAI21_X1 _31169_ (.A(_07582_),
    .B1(_07583_),
    .B2(_07584_),
    .ZN(_07585_));
 AOI221_X2 _31170_ (.A(_19626_),
    .B1(_07535_),
    .B2(_07585_),
    .C1(_07522_),
    .C2(_19628_),
    .ZN(_07586_));
 XNOR2_X2 _31171_ (.A(_07508_),
    .B(_07586_),
    .ZN(_07587_));
 XNOR2_X1 _31172_ (.A(_07514_),
    .B(_07585_),
    .ZN(_07588_));
 NOR3_X1 _31173_ (.A1(_07494_),
    .A2(_07499_),
    .A3(_07588_),
    .ZN(_07589_));
 XNOR2_X2 _31174_ (.A(_07522_),
    .B(_07579_),
    .ZN(_07590_));
 AND3_X1 _31175_ (.A1(_07587_),
    .A2(_07589_),
    .A3(_07590_),
    .ZN(_07591_));
 NAND2_X1 _31176_ (.A1(_07508_),
    .A2(_07522_),
    .ZN(_07592_));
 OAI21_X1 _31177_ (.A(_07509_),
    .B1(_07515_),
    .B2(_07592_),
    .ZN(_07593_));
 NOR2_X1 _31178_ (.A1(_07577_),
    .A2(_07592_),
    .ZN(_07594_));
 AOI21_X2 _31179_ (.A(_07593_),
    .B1(_07594_),
    .B2(_07493_),
    .ZN(_07595_));
 XNOR2_X2 _31180_ (.A(_07510_),
    .B(_07595_),
    .ZN(_07596_));
 INV_X1 _31181_ (.A(_07506_),
    .ZN(_07597_));
 NAND4_X1 _31182_ (.A1(_07510_),
    .A2(_07508_),
    .A3(_07535_),
    .A4(_07585_),
    .ZN(_07598_));
 NAND2_X1 _31183_ (.A1(_07534_),
    .A2(_07598_),
    .ZN(_07599_));
 XNOR2_X1 _31184_ (.A(_07597_),
    .B(_07599_),
    .ZN(_07600_));
 NAND3_X1 _31185_ (.A1(_07591_),
    .A2(_07596_),
    .A3(_07600_),
    .ZN(_07601_));
 OR3_X1 _31186_ (.A1(_07576_),
    .A2(_07581_),
    .A3(_07601_),
    .ZN(_07602_));
 INV_X1 _31187_ (.A(_07504_),
    .ZN(_07603_));
 NOR3_X1 _31188_ (.A1(_07517_),
    .A2(_07467_),
    .A3(_07469_),
    .ZN(_07604_));
 AOI21_X1 _31189_ (.A(_07452_),
    .B1(_19646_),
    .B2(_07457_),
    .ZN(_07605_));
 OAI21_X1 _31190_ (.A(_07470_),
    .B1(_07475_),
    .B2(_07605_),
    .ZN(_07606_));
 AOI221_X2 _31191_ (.A(_19632_),
    .B1(_07488_),
    .B2(_07490_),
    .C1(_07604_),
    .C2(_07606_),
    .ZN(_07607_));
 NOR3_X1 _31192_ (.A1(_07577_),
    .A2(_07592_),
    .A3(_07607_),
    .ZN(_07608_));
 OAI21_X1 _31193_ (.A(_07510_),
    .B1(_07593_),
    .B2(_07608_),
    .ZN(_07609_));
 AOI21_X1 _31194_ (.A(_07597_),
    .B1(_07507_),
    .B2(_07609_),
    .ZN(_07610_));
 OAI21_X1 _31195_ (.A(_07525_),
    .B1(_07610_),
    .B2(_07505_),
    .ZN(_07611_));
 AOI21_X1 _31196_ (.A(_07503_),
    .B1(_07603_),
    .B2(_07611_),
    .ZN(_07612_));
 NOR2_X1 _31197_ (.A1(_19616_),
    .A2(_07612_),
    .ZN(_07613_));
 XNOR2_X2 _31198_ (.A(_19615_),
    .B(_07613_),
    .ZN(_07614_));
 INV_X1 _31199_ (.A(_07614_),
    .ZN(_07615_));
 NOR2_X1 _31200_ (.A1(_07602_),
    .A2(_07615_),
    .ZN(_07616_));
 NAND2_X1 _31201_ (.A1(_07553_),
    .A2(_07616_),
    .ZN(_07617_));
 XNOR2_X1 _31202_ (.A(_07529_),
    .B(_07617_),
    .ZN(_14275_));
 INV_X1 _31203_ (.A(_14275_),
    .ZN(_14280_));
 INV_X2 _31204_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.b ),
    .ZN(_07618_));
 CLKBUF_X3 _31205_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.b ),
    .Z(_07619_));
 NOR4_X2 _31206_ (.A1(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07619_),
    .ZN(_07620_));
 NAND2_X4 _31207_ (.A1(_07618_),
    .A2(_07620_),
    .ZN(_07621_));
 OR4_X1 _31208_ (.A1(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07622_));
 OAI21_X2 _31209_ (.A(_07621_),
    .B1(_07622_),
    .B2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07623_));
 NAND4_X2 _31210_ (.A1(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.b ),
    .A2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .A3(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .A4(_07619_),
    .ZN(_07624_));
 NOR2_X4 _31211_ (.A1(_07618_),
    .A2(_07624_),
    .ZN(_07625_));
 AND4_X1 _31212_ (.A1(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07626_));
 AOI21_X4 _31213_ (.A(_07625_),
    .B1(_07626_),
    .B2(\g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07627_));
 INV_X1 _31214_ (.A(_14277_),
    .ZN(_07628_));
 AOI21_X1 _31215_ (.A(_07623_),
    .B1(_07627_),
    .B2(_07628_),
    .ZN(_00241_));
 INV_X1 _31216_ (.A(_19655_),
    .ZN(_07629_));
 AOI21_X1 _31217_ (.A(_07623_),
    .B1(_07627_),
    .B2(_07629_),
    .ZN(_00242_));
 INV_X1 _31218_ (.A(_14286_),
    .ZN(_07630_));
 AOI21_X1 _31219_ (.A(_07623_),
    .B1(_07627_),
    .B2(_07630_),
    .ZN(_00243_));
 XOR2_X1 _31220_ (.A(_14285_),
    .B(_19664_),
    .Z(_07631_));
 AOI21_X1 _31221_ (.A(_07623_),
    .B1(_07627_),
    .B2(_07631_),
    .ZN(_00244_));
 AOI21_X1 _31222_ (.A(_19659_),
    .B1(_19660_),
    .B2(_19654_),
    .ZN(_07632_));
 INV_X1 _31223_ (.A(_07632_),
    .ZN(_07633_));
 AOI21_X1 _31224_ (.A(_19663_),
    .B1(_07633_),
    .B2(_19664_),
    .ZN(_07634_));
 XNOR2_X1 _31225_ (.A(_07619_),
    .B(_19661_),
    .ZN(_07635_));
 XNOR2_X1 _31226_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_07635_),
    .ZN(_07636_));
 XNOR2_X1 _31227_ (.A(_07634_),
    .B(_07636_),
    .ZN(_07637_));
 AOI21_X1 _31228_ (.A(_07623_),
    .B1(_07627_),
    .B2(_07637_),
    .ZN(_00245_));
 INV_X1 _31229_ (.A(_07623_),
    .ZN(_07638_));
 NAND2_X4 _31230_ (.A1(_07638_),
    .A2(_07627_),
    .ZN(_07639_));
 INV_X1 _31231_ (.A(_07639_),
    .ZN(_07640_));
 NAND2_X1 _31232_ (.A1(_07496_),
    .A2(_07640_),
    .ZN(_07641_));
 NOR2_X1 _31233_ (.A1(_07499_),
    .A2(_07641_),
    .ZN(_07642_));
 AND2_X1 _31234_ (.A1(_19668_),
    .A2(_07640_),
    .ZN(_07643_));
 MUX2_X1 _31235_ (.A(_07642_),
    .B(_07643_),
    .S(_14275_),
    .Z(_00240_));
 XOR2_X1 _31236_ (.A(_19667_),
    .B(_07588_),
    .Z(_07644_));
 NOR2_X1 _31237_ (.A1(_07639_),
    .A2(_07644_),
    .ZN(_07645_));
 MUX2_X1 _31238_ (.A(_07643_),
    .B(_07645_),
    .S(_14275_),
    .Z(_00246_));
 XNOR2_X1 _31239_ (.A(_07589_),
    .B(_07590_),
    .ZN(_07646_));
 NOR2_X1 _31240_ (.A1(_07639_),
    .A2(_07646_),
    .ZN(_07647_));
 MUX2_X1 _31241_ (.A(_07645_),
    .B(_07647_),
    .S(_14275_),
    .Z(_00247_));
 NAND2_X1 _31242_ (.A1(_19667_),
    .A2(_07590_),
    .ZN(_07648_));
 NOR2_X1 _31243_ (.A1(_07588_),
    .A2(_07648_),
    .ZN(_07649_));
 XNOR2_X1 _31244_ (.A(_07587_),
    .B(_07649_),
    .ZN(_07650_));
 NOR2_X1 _31245_ (.A1(_07639_),
    .A2(_07650_),
    .ZN(_07651_));
 MUX2_X1 _31246_ (.A(_07647_),
    .B(_07651_),
    .S(_14275_),
    .Z(_00248_));
 XNOR2_X1 _31247_ (.A(_07591_),
    .B(_07596_),
    .ZN(_07652_));
 NOR2_X1 _31248_ (.A1(_07639_),
    .A2(_07652_),
    .ZN(_07653_));
 MUX2_X1 _31249_ (.A(_07651_),
    .B(_07653_),
    .S(_14275_),
    .Z(_00249_));
 INV_X1 _31250_ (.A(_07600_),
    .ZN(_07654_));
 NAND3_X1 _31251_ (.A1(_07587_),
    .A2(_07596_),
    .A3(_07649_),
    .ZN(_07655_));
 XNOR2_X1 _31252_ (.A(_07654_),
    .B(_07655_),
    .ZN(_07656_));
 NOR2_X1 _31253_ (.A1(_07639_),
    .A2(_07656_),
    .ZN(_07657_));
 MUX2_X1 _31254_ (.A(_07653_),
    .B(_07657_),
    .S(_14275_),
    .Z(_00250_));
 XNOR2_X1 _31255_ (.A(_07581_),
    .B(_07601_),
    .ZN(_07658_));
 NOR2_X1 _31256_ (.A1(_07639_),
    .A2(_07658_),
    .ZN(_07659_));
 MUX2_X1 _31257_ (.A(_07657_),
    .B(_07659_),
    .S(_14275_),
    .Z(_00251_));
 OR3_X2 _31258_ (.A1(_07581_),
    .A2(_07654_),
    .A3(_07655_),
    .ZN(_07660_));
 XNOR2_X2 _31259_ (.A(_07576_),
    .B(_07660_),
    .ZN(_07661_));
 NOR2_X1 _31260_ (.A1(_07639_),
    .A2(_07661_),
    .ZN(_07662_));
 MUX2_X1 _31261_ (.A(_07659_),
    .B(_07662_),
    .S(_14275_),
    .Z(_00252_));
 AOI21_X1 _31262_ (.A(_07639_),
    .B1(_07661_),
    .B2(_07616_),
    .ZN(_07663_));
 AOI21_X1 _31263_ (.A(_07661_),
    .B1(_07616_),
    .B2(_07553_),
    .ZN(_07664_));
 INV_X1 _31264_ (.A(_07602_),
    .ZN(_07665_));
 NOR2_X1 _31265_ (.A1(_07665_),
    .A2(_07614_),
    .ZN(_07666_));
 INV_X1 _31266_ (.A(_07553_),
    .ZN(_07667_));
 AOI21_X1 _31267_ (.A(_07666_),
    .B1(_07616_),
    .B2(_07667_),
    .ZN(_07668_));
 MUX2_X1 _31268_ (.A(_07664_),
    .B(_07668_),
    .S(_07529_),
    .Z(_07669_));
 AND2_X1 _31269_ (.A1(_07663_),
    .A2(_07669_),
    .ZN(_00253_));
 OAI21_X1 _31270_ (.A(_07553_),
    .B1(_07660_),
    .B2(_07576_),
    .ZN(_07670_));
 AOI21_X1 _31271_ (.A(_07666_),
    .B1(_07670_),
    .B2(_07616_),
    .ZN(_07671_));
 NOR2_X1 _31272_ (.A1(_07576_),
    .A2(_07660_),
    .ZN(_07672_));
 OAI21_X1 _31273_ (.A(_07614_),
    .B1(_07672_),
    .B2(_07665_),
    .ZN(_07673_));
 NOR3_X1 _31274_ (.A1(_07576_),
    .A2(_07615_),
    .A3(_07660_),
    .ZN(_07674_));
 MUX2_X1 _31275_ (.A(_07673_),
    .B(_07674_),
    .S(_07667_),
    .Z(_07675_));
 MUX2_X1 _31276_ (.A(_07671_),
    .B(_07675_),
    .S(_07529_),
    .Z(_07676_));
 AND2_X1 _31277_ (.A1(_07640_),
    .A2(_07676_),
    .ZN(_00254_));
 CLKBUF_X2 _31278_ (.A(_19692_),
    .Z(_07677_));
 AOI21_X1 _31279_ (.A(_19691_),
    .B1(_07677_),
    .B2(_19693_),
    .ZN(_07678_));
 BUF_X1 _31280_ (.A(_19694_),
    .Z(_07679_));
 NAND2_X1 _31281_ (.A1(_07677_),
    .A2(_07679_),
    .ZN(_07680_));
 CLKBUF_X2 _31282_ (.A(_19697_),
    .Z(_07681_));
 AOI21_X1 _31283_ (.A(_19695_),
    .B1(_19696_),
    .B2(_07681_),
    .ZN(_07682_));
 OAI21_X1 _31284_ (.A(_07678_),
    .B1(_07680_),
    .B2(_07682_),
    .ZN(_07683_));
 INV_X1 _31285_ (.A(_19699_),
    .ZN(_07684_));
 CLKBUF_X2 _31286_ (.A(_19701_),
    .Z(_07685_));
 INV_X1 _31287_ (.A(_19703_),
    .ZN(_07686_));
 AOI21_X1 _31288_ (.A(_19705_),
    .B1(_19706_),
    .B2(_19707_),
    .ZN(_07687_));
 INV_X1 _31289_ (.A(_19704_),
    .ZN(_07688_));
 OAI21_X1 _31290_ (.A(_07686_),
    .B1(_07687_),
    .B2(_07688_),
    .ZN(_07689_));
 CLKBUF_X2 _31291_ (.A(_19702_),
    .Z(_07690_));
 AOI21_X1 _31292_ (.A(_07685_),
    .B1(_07689_),
    .B2(_07690_),
    .ZN(_07691_));
 INV_X1 _31293_ (.A(_19700_),
    .ZN(_07692_));
 OAI21_X2 _31294_ (.A(_07684_),
    .B1(_07691_),
    .B2(_07692_),
    .ZN(_07693_));
 INV_X1 _31295_ (.A(_19696_),
    .ZN(_07694_));
 BUF_X2 _31296_ (.A(_19698_),
    .Z(_07695_));
 INV_X1 _31297_ (.A(_07695_),
    .ZN(_07696_));
 NOR3_X2 _31298_ (.A1(_07694_),
    .A2(_07696_),
    .A3(_07680_),
    .ZN(_07697_));
 AOI21_X2 _31299_ (.A(_07683_),
    .B1(_07693_),
    .B2(_07697_),
    .ZN(_07698_));
 XNOR2_X1 _31300_ (.A(_19690_),
    .B(_07698_),
    .ZN(_07699_));
 INV_X1 _31301_ (.A(_19695_),
    .ZN(_07700_));
 AOI21_X1 _31302_ (.A(_07681_),
    .B1(_07695_),
    .B2(_07693_),
    .ZN(_07701_));
 OAI21_X2 _31303_ (.A(_07700_),
    .B1(_07701_),
    .B2(_07694_),
    .ZN(_07702_));
 XNOR2_X1 _31304_ (.A(_07679_),
    .B(_07702_),
    .ZN(_07703_));
 XNOR2_X1 _31305_ (.A(_07695_),
    .B(_07693_),
    .ZN(_07704_));
 INV_X1 _31306_ (.A(_19689_),
    .ZN(_07705_));
 INV_X1 _31307_ (.A(_19690_),
    .ZN(_07706_));
 AOI21_X1 _31308_ (.A(_19693_),
    .B1(_07679_),
    .B2(_19695_),
    .ZN(_07707_));
 INV_X1 _31309_ (.A(_07707_),
    .ZN(_07708_));
 AOI21_X1 _31310_ (.A(_19691_),
    .B1(_07708_),
    .B2(_07677_),
    .ZN(_07709_));
 OAI21_X1 _31311_ (.A(_07705_),
    .B1(_07706_),
    .B2(_07709_),
    .ZN(_07710_));
 INV_X1 _31312_ (.A(_07677_),
    .ZN(_07711_));
 NAND2_X1 _31313_ (.A1(_07679_),
    .A2(_19696_),
    .ZN(_07712_));
 NOR3_X2 _31314_ (.A1(_07706_),
    .A2(_07711_),
    .A3(_07712_),
    .ZN(_07713_));
 AOI21_X2 _31315_ (.A(_07681_),
    .B1(_07695_),
    .B2(_19699_),
    .ZN(_07714_));
 OAI21_X1 _31316_ (.A(_07686_),
    .B1(_07688_),
    .B2(_14290_),
    .ZN(_07715_));
 AOI21_X1 _31317_ (.A(_07685_),
    .B1(_07715_),
    .B2(_07690_),
    .ZN(_07716_));
 NAND2_X1 _31318_ (.A1(_07695_),
    .A2(_19700_),
    .ZN(_07717_));
 NOR2_X1 _31319_ (.A1(_07716_),
    .A2(_07717_),
    .ZN(_07718_));
 INV_X1 _31320_ (.A(_07718_),
    .ZN(_07719_));
 NAND2_X1 _31321_ (.A1(_07714_),
    .A2(_07719_),
    .ZN(_07720_));
 AOI21_X1 _31322_ (.A(_07710_),
    .B1(_07713_),
    .B2(_07720_),
    .ZN(_07721_));
 XNOR2_X1 _31323_ (.A(_19688_),
    .B(_07721_),
    .ZN(_19722_));
 AOI21_X1 _31324_ (.A(_07696_),
    .B1(_07692_),
    .B2(_07684_),
    .ZN(_07722_));
 NOR2_X1 _31325_ (.A1(_07681_),
    .A2(_07722_),
    .ZN(_07723_));
 XNOR2_X1 _31326_ (.A(_07694_),
    .B(_07723_),
    .ZN(_07724_));
 XNOR2_X1 _31327_ (.A(_14290_),
    .B(_19704_),
    .ZN(_07725_));
 NOR4_X1 _31328_ (.A1(_14291_),
    .A2(\g_row[1].g_col[0].mult.adder.a[0] ),
    .A3(_19708_),
    .A4(_07725_),
    .ZN(_07726_));
 XNOR2_X1 _31329_ (.A(_07692_),
    .B(_07716_),
    .ZN(_07727_));
 XNOR2_X1 _31330_ (.A(_07690_),
    .B(_07689_),
    .ZN(_07728_));
 NAND4_X1 _31331_ (.A1(_07724_),
    .A2(_07726_),
    .A3(_07727_),
    .A4(_07728_),
    .ZN(_07729_));
 OAI21_X1 _31332_ (.A(_07707_),
    .B1(_07712_),
    .B2(_07714_),
    .ZN(_07730_));
 NOR2_X1 _31333_ (.A1(_07712_),
    .A2(_07719_),
    .ZN(_07731_));
 NOR2_X1 _31334_ (.A1(_07730_),
    .A2(_07731_),
    .ZN(_07732_));
 XNOR2_X1 _31335_ (.A(_07677_),
    .B(_07732_),
    .ZN(_07733_));
 NOR3_X1 _31336_ (.A1(_19722_),
    .A2(_07729_),
    .A3(_07733_),
    .ZN(_07734_));
 NAND3_X1 _31337_ (.A1(_07703_),
    .A2(_07704_),
    .A3(_07734_),
    .ZN(_07735_));
 AND2_X1 _31338_ (.A1(_07699_),
    .A2(_07735_),
    .ZN(_19723_));
 INV_X1 _31339_ (.A(_19669_),
    .ZN(_07736_));
 INV_X1 _31340_ (.A(_19670_),
    .ZN(_07737_));
 INV_X1 _31341_ (.A(_19673_),
    .ZN(_07738_));
 INV_X1 _31342_ (.A(_19674_),
    .ZN(_07739_));
 INV_X1 _31343_ (.A(_19679_),
    .ZN(_07740_));
 BUF_X2 _31344_ (.A(_19682_),
    .Z(_07741_));
 AOI21_X2 _31345_ (.A(_19681_),
    .B1(_07741_),
    .B2(_19683_),
    .ZN(_07742_));
 CLKBUF_X2 _31346_ (.A(_19680_),
    .Z(_07743_));
 INV_X1 _31347_ (.A(_07743_),
    .ZN(_07744_));
 OAI21_X1 _31348_ (.A(_07740_),
    .B1(_07742_),
    .B2(_07744_),
    .ZN(_07745_));
 AOI21_X1 _31349_ (.A(_19677_),
    .B1(_19678_),
    .B2(_07745_),
    .ZN(_07746_));
 BUF_X2 _31350_ (.A(_19686_),
    .Z(_07747_));
 AND2_X1 _31351_ (.A1(_07747_),
    .A2(_19688_),
    .ZN(_07748_));
 AOI21_X1 _31352_ (.A(_19691_),
    .B1(_07730_),
    .B2(_07677_),
    .ZN(_07749_));
 OAI21_X1 _31353_ (.A(_07705_),
    .B1(_07706_),
    .B2(_07749_),
    .ZN(_07750_));
 AOI221_X2 _31354_ (.A(_19685_),
    .B1(_07747_),
    .B2(_19687_),
    .C1(_07748_),
    .C2(_07750_),
    .ZN(_07751_));
 BUF_X2 _31355_ (.A(_19684_),
    .Z(_07752_));
 NAND4_X1 _31356_ (.A1(_19678_),
    .A2(_07743_),
    .A3(_07741_),
    .A4(_07752_),
    .ZN(_07753_));
 OAI21_X1 _31357_ (.A(_07746_),
    .B1(_07751_),
    .B2(_07753_),
    .ZN(_07754_));
 BUF_X2 _31358_ (.A(_19676_),
    .Z(_07755_));
 AOI21_X1 _31359_ (.A(_19675_),
    .B1(_07754_),
    .B2(_07755_),
    .ZN(_07756_));
 OAI21_X1 _31360_ (.A(_07738_),
    .B1(_07739_),
    .B2(_07756_),
    .ZN(_07757_));
 AOI21_X1 _31361_ (.A(_19671_),
    .B1(_19672_),
    .B2(_07757_),
    .ZN(_07758_));
 OAI21_X2 _31362_ (.A(_07736_),
    .B1(_07737_),
    .B2(_07758_),
    .ZN(_07759_));
 INV_X1 _31363_ (.A(_19681_),
    .ZN(_07760_));
 INV_X1 _31364_ (.A(_07741_),
    .ZN(_07761_));
 AOI21_X1 _31365_ (.A(_19683_),
    .B1(_07752_),
    .B2(_19685_),
    .ZN(_07762_));
 OAI21_X1 _31366_ (.A(_07760_),
    .B1(_07761_),
    .B2(_07762_),
    .ZN(_07763_));
 AOI21_X1 _31367_ (.A(_19679_),
    .B1(_07763_),
    .B2(_07743_),
    .ZN(_07764_));
 NAND4_X1 _31368_ (.A1(_07743_),
    .A2(_07741_),
    .A3(_07752_),
    .A4(_07747_),
    .ZN(_07765_));
 AOI21_X1 _31369_ (.A(_19687_),
    .B1(_19688_),
    .B2(_19689_),
    .ZN(_07766_));
 NAND2_X1 _31370_ (.A1(_19688_),
    .A2(_19690_),
    .ZN(_07767_));
 OAI21_X1 _31371_ (.A(_07766_),
    .B1(_07767_),
    .B2(_07678_),
    .ZN(_07768_));
 NOR2_X1 _31372_ (.A1(_07680_),
    .A2(_07767_),
    .ZN(_07769_));
 INV_X1 _31373_ (.A(_07685_),
    .ZN(_07770_));
 OAI21_X1 _31374_ (.A(_07684_),
    .B1(_07770_),
    .B2(_07692_),
    .ZN(_07771_));
 AOI21_X1 _31375_ (.A(_07681_),
    .B1(_07695_),
    .B2(_07771_),
    .ZN(_07772_));
 OAI21_X1 _31376_ (.A(_07700_),
    .B1(_07772_),
    .B2(_07694_),
    .ZN(_07773_));
 AOI21_X1 _31377_ (.A(_07768_),
    .B1(_07769_),
    .B2(_07773_),
    .ZN(_07774_));
 OAI21_X1 _31378_ (.A(_07764_),
    .B1(_07765_),
    .B2(_07774_),
    .ZN(_07775_));
 AOI21_X1 _31379_ (.A(_19677_),
    .B1(_19678_),
    .B2(_07775_),
    .ZN(_07776_));
 INV_X1 _31380_ (.A(_07776_),
    .ZN(_07777_));
 AOI21_X1 _31381_ (.A(_19675_),
    .B1(_07777_),
    .B2(_07755_),
    .ZN(_07778_));
 OAI21_X1 _31382_ (.A(_07738_),
    .B1(_07739_),
    .B2(_07778_),
    .ZN(_07779_));
 AOI21_X2 _31383_ (.A(_19671_),
    .B1(_19672_),
    .B2(_07779_),
    .ZN(_07780_));
 XNOR2_X2 _31384_ (.A(_19670_),
    .B(_07780_),
    .ZN(_07781_));
 NAND2_X1 _31385_ (.A1(_07713_),
    .A2(_07748_),
    .ZN(_07782_));
 OAI21_X2 _31386_ (.A(_07751_),
    .B1(_07782_),
    .B2(_07719_),
    .ZN(_07783_));
 INV_X1 _31387_ (.A(_07783_),
    .ZN(_07784_));
 OAI21_X1 _31388_ (.A(_07746_),
    .B1(_07753_),
    .B2(_07784_),
    .ZN(_07785_));
 XOR2_X2 _31389_ (.A(_07755_),
    .B(_07785_),
    .Z(_07786_));
 INV_X1 _31390_ (.A(_19677_),
    .ZN(_07787_));
 INV_X1 _31391_ (.A(_19678_),
    .ZN(_07788_));
 NAND2_X1 _31392_ (.A1(_07752_),
    .A2(_07747_),
    .ZN(_07789_));
 OAI21_X1 _31393_ (.A(_07762_),
    .B1(_07789_),
    .B2(_07766_),
    .ZN(_07790_));
 INV_X1 _31394_ (.A(_19705_),
    .ZN(_07791_));
 OAI21_X1 _31395_ (.A(_07686_),
    .B1(_07791_),
    .B2(_07688_),
    .ZN(_07792_));
 AOI21_X1 _31396_ (.A(_07685_),
    .B1(_07792_),
    .B2(_07690_),
    .ZN(_07793_));
 OAI21_X1 _31397_ (.A(_07684_),
    .B1(_07793_),
    .B2(_07692_),
    .ZN(_07794_));
 AOI21_X1 _31398_ (.A(_07683_),
    .B1(_07697_),
    .B2(_07794_),
    .ZN(_07795_));
 NOR3_X1 _31399_ (.A1(_07789_),
    .A2(_07767_),
    .A3(_07795_),
    .ZN(_07796_));
 OAI21_X1 _31400_ (.A(_07741_),
    .B1(_07790_),
    .B2(_07796_),
    .ZN(_07797_));
 NAND2_X1 _31401_ (.A1(_07760_),
    .A2(_07797_),
    .ZN(_07798_));
 AOI21_X1 _31402_ (.A(_19679_),
    .B1(_07798_),
    .B2(_07743_),
    .ZN(_07799_));
 OAI21_X1 _31403_ (.A(_07787_),
    .B1(_07788_),
    .B2(_07799_),
    .ZN(_07800_));
 AOI21_X2 _31404_ (.A(_19675_),
    .B1(_07800_),
    .B2(_07755_),
    .ZN(_07801_));
 XNOR2_X2 _31405_ (.A(_19674_),
    .B(_07801_),
    .ZN(_07802_));
 AOI21_X2 _31406_ (.A(_19685_),
    .B1(_07747_),
    .B2(_19687_),
    .ZN(_07803_));
 NAND2_X1 _31407_ (.A1(_07741_),
    .A2(_07752_),
    .ZN(_07804_));
 NAND3_X1 _31408_ (.A1(_07741_),
    .A2(_07752_),
    .A3(_07748_),
    .ZN(_07805_));
 OAI221_X2 _31409_ (.A(_07742_),
    .B1(_07803_),
    .B2(_07804_),
    .C1(_07805_),
    .C2(_07721_),
    .ZN(_07806_));
 XNOR2_X2 _31410_ (.A(_07744_),
    .B(_07806_),
    .ZN(_07807_));
 AOI21_X2 _31411_ (.A(_07768_),
    .B1(_07769_),
    .B2(_07702_),
    .ZN(_07808_));
 XNOR2_X2 _31412_ (.A(_07747_),
    .B(_07808_),
    .ZN(_07809_));
 AND3_X1 _31413_ (.A1(_07699_),
    .A2(_19722_),
    .A3(_07809_),
    .ZN(_07810_));
 NOR3_X1 _31414_ (.A1(_07698_),
    .A2(_07789_),
    .A3(_07767_),
    .ZN(_07811_));
 NOR2_X1 _31415_ (.A1(_07790_),
    .A2(_07811_),
    .ZN(_07812_));
 XNOR2_X2 _31416_ (.A(_07761_),
    .B(_07812_),
    .ZN(_07813_));
 INV_X1 _31417_ (.A(_07813_),
    .ZN(_07814_));
 XOR2_X2 _31418_ (.A(_07752_),
    .B(_07783_),
    .Z(_07815_));
 AND3_X1 _31419_ (.A1(_07810_),
    .A2(_07814_),
    .A3(_07815_),
    .ZN(_07816_));
 OAI21_X1 _31420_ (.A(_07764_),
    .B1(_07765_),
    .B2(_07808_),
    .ZN(_07817_));
 XNOR2_X2 _31421_ (.A(_07788_),
    .B(_07817_),
    .ZN(_07818_));
 NAND3_X1 _31422_ (.A1(_07807_),
    .A2(_07816_),
    .A3(_07818_),
    .ZN(_07819_));
 INV_X1 _31423_ (.A(_07819_),
    .ZN(_07820_));
 NAND3_X1 _31424_ (.A1(_07786_),
    .A2(_07802_),
    .A3(_07820_),
    .ZN(_07821_));
 AOI21_X1 _31425_ (.A(_07685_),
    .B1(_19703_),
    .B2(_07690_),
    .ZN(_07822_));
 OAI21_X1 _31426_ (.A(_07714_),
    .B1(_07717_),
    .B2(_07822_),
    .ZN(_07823_));
 AOI21_X1 _31427_ (.A(_07710_),
    .B1(_07713_),
    .B2(_07823_),
    .ZN(_07824_));
 OAI221_X1 _31428_ (.A(_07742_),
    .B1(_07803_),
    .B2(_07804_),
    .C1(_07805_),
    .C2(_07824_),
    .ZN(_07825_));
 AOI21_X1 _31429_ (.A(_19679_),
    .B1(_07825_),
    .B2(_07743_),
    .ZN(_07826_));
 OAI21_X1 _31430_ (.A(_07787_),
    .B1(_07788_),
    .B2(_07826_),
    .ZN(_07827_));
 AOI21_X1 _31431_ (.A(_19675_),
    .B1(_07827_),
    .B2(_07755_),
    .ZN(_07828_));
 OAI21_X1 _31432_ (.A(_07738_),
    .B1(_07739_),
    .B2(_07828_),
    .ZN(_07829_));
 XNOR2_X2 _31433_ (.A(_19672_),
    .B(_07829_),
    .ZN(_07830_));
 OR2_X1 _31434_ (.A1(_07821_),
    .A2(_07830_),
    .ZN(_07831_));
 INV_X1 _31435_ (.A(_07831_),
    .ZN(_07832_));
 NAND2_X1 _31436_ (.A1(_07781_),
    .A2(_07832_),
    .ZN(_07833_));
 XNOR2_X1 _31437_ (.A(_07759_),
    .B(_07833_),
    .ZN(_07834_));
 BUF_X1 _31438_ (.A(_07834_),
    .Z(_14293_));
 INV_X1 _31439_ (.A(_14293_),
    .ZN(_14297_));
 OR4_X1 _31440_ (.A1(\g_row[1].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07835_));
 OAI21_X2 _31441_ (.A(_06947_),
    .B1(_07835_),
    .B2(\g_row[1].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07836_));
 AND4_X1 _31442_ (.A1(\g_row[1].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_07837_));
 AOI21_X4 _31443_ (.A(_06951_),
    .B1(_07837_),
    .B2(\g_row[1].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_07838_));
 INV_X1 _31444_ (.A(_14295_),
    .ZN(_07839_));
 AOI21_X1 _31445_ (.A(_07836_),
    .B1(_07838_),
    .B2(_07839_),
    .ZN(_00257_));
 INV_X1 _31446_ (.A(_19712_),
    .ZN(_07840_));
 AOI21_X1 _31447_ (.A(_07836_),
    .B1(_07838_),
    .B2(_07840_),
    .ZN(_00258_));
 INV_X1 _31448_ (.A(_14303_),
    .ZN(_07841_));
 AOI21_X1 _31449_ (.A(_07836_),
    .B1(_07838_),
    .B2(_07841_),
    .ZN(_00259_));
 XOR2_X1 _31450_ (.A(_14302_),
    .B(_19721_),
    .Z(_07842_));
 AOI21_X1 _31451_ (.A(_07836_),
    .B1(_07838_),
    .B2(_07842_),
    .ZN(_00260_));
 AOI21_X1 _31452_ (.A(_19716_),
    .B1(_19717_),
    .B2(_19711_),
    .ZN(_07843_));
 INV_X1 _31453_ (.A(_07843_),
    .ZN(_07844_));
 AOI21_X1 _31454_ (.A(_19720_),
    .B1(_07844_),
    .B2(_19721_),
    .ZN(_07845_));
 XNOR2_X1 _31455_ (.A(\g_row[1].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_19718_),
    .ZN(_07846_));
 XNOR2_X1 _31456_ (.A(_06945_),
    .B(_07846_),
    .ZN(_07847_));
 XNOR2_X1 _31457_ (.A(_07845_),
    .B(_07847_),
    .ZN(_07848_));
 AOI21_X1 _31458_ (.A(_07836_),
    .B1(_07838_),
    .B2(_07848_),
    .ZN(_00261_));
 INV_X1 _31459_ (.A(_07836_),
    .ZN(_07849_));
 NAND2_X4 _31460_ (.A1(_07849_),
    .A2(_07838_),
    .ZN(_07850_));
 INV_X1 _31461_ (.A(_07699_),
    .ZN(_07851_));
 NOR3_X1 _31462_ (.A1(_07851_),
    .A2(_07735_),
    .A3(_07834_),
    .ZN(_07852_));
 AOI21_X1 _31463_ (.A(_07852_),
    .B1(_14293_),
    .B2(_19725_),
    .ZN(_07853_));
 NOR2_X1 _31464_ (.A1(_07850_),
    .A2(_07853_),
    .ZN(_00256_));
 XNOR2_X1 _31465_ (.A(_19724_),
    .B(_07809_),
    .ZN(_07854_));
 NAND2_X1 _31466_ (.A1(_14293_),
    .A2(_07854_),
    .ZN(_07855_));
 OAI21_X2 _31467_ (.A(_07855_),
    .B1(_14293_),
    .B2(_19725_),
    .ZN(_07856_));
 NOR2_X1 _31468_ (.A1(_07850_),
    .A2(_07856_),
    .ZN(_00262_));
 XNOR2_X1 _31469_ (.A(_07810_),
    .B(_07815_),
    .ZN(_07857_));
 MUX2_X1 _31470_ (.A(_07854_),
    .B(_07857_),
    .S(_14293_),
    .Z(_07858_));
 NOR2_X1 _31471_ (.A1(_07850_),
    .A2(_07858_),
    .ZN(_00263_));
 NAND3_X1 _31472_ (.A1(_19724_),
    .A2(_07809_),
    .A3(_07815_),
    .ZN(_07859_));
 XNOR2_X1 _31473_ (.A(_07813_),
    .B(_07859_),
    .ZN(_07860_));
 MUX2_X1 _31474_ (.A(_07857_),
    .B(_07860_),
    .S(_14293_),
    .Z(_07861_));
 NOR2_X1 _31475_ (.A1(_07850_),
    .A2(_07861_),
    .ZN(_00264_));
 XNOR2_X1 _31476_ (.A(_07807_),
    .B(_07816_),
    .ZN(_07862_));
 MUX2_X1 _31477_ (.A(_07860_),
    .B(_07862_),
    .S(_14293_),
    .Z(_07863_));
 NOR2_X1 _31478_ (.A1(_07850_),
    .A2(_07863_),
    .ZN(_00265_));
 INV_X1 _31479_ (.A(_07807_),
    .ZN(_07864_));
 NOR3_X1 _31480_ (.A1(_07864_),
    .A2(_07813_),
    .A3(_07859_),
    .ZN(_07865_));
 XNOR2_X1 _31481_ (.A(_07818_),
    .B(_07865_),
    .ZN(_07866_));
 MUX2_X1 _31482_ (.A(_07862_),
    .B(_07866_),
    .S(_07834_),
    .Z(_07867_));
 NOR2_X1 _31483_ (.A1(_07850_),
    .A2(_07867_),
    .ZN(_00266_));
 XOR2_X1 _31484_ (.A(_07786_),
    .B(_07819_),
    .Z(_07868_));
 MUX2_X1 _31485_ (.A(_07866_),
    .B(_07868_),
    .S(_07834_),
    .Z(_07869_));
 NOR2_X1 _31486_ (.A1(_07850_),
    .A2(_07869_),
    .ZN(_00267_));
 NOR2_X1 _31487_ (.A1(_14293_),
    .A2(_07868_),
    .ZN(_07870_));
 NAND3_X1 _31488_ (.A1(_07786_),
    .A2(_07818_),
    .A3(_07865_),
    .ZN(_07871_));
 XNOR2_X2 _31489_ (.A(_07802_),
    .B(_07871_),
    .ZN(_07872_));
 AOI21_X2 _31490_ (.A(_07870_),
    .B1(_07872_),
    .B2(_14293_),
    .ZN(_07873_));
 NOR2_X1 _31491_ (.A1(_07850_),
    .A2(_07873_),
    .ZN(_00268_));
 NOR2_X1 _31492_ (.A1(_07831_),
    .A2(_07872_),
    .ZN(_07874_));
 NAND2_X1 _31493_ (.A1(_07833_),
    .A2(_07872_),
    .ZN(_07875_));
 NAND2_X1 _31494_ (.A1(_07821_),
    .A2(_07830_),
    .ZN(_07876_));
 OAI21_X1 _31495_ (.A(_07876_),
    .B1(_07831_),
    .B2(_07781_),
    .ZN(_07877_));
 MUX2_X1 _31496_ (.A(_07875_),
    .B(_07877_),
    .S(_07759_),
    .Z(_07878_));
 NOR3_X1 _31497_ (.A1(_07850_),
    .A2(_07874_),
    .A3(_07878_),
    .ZN(_00269_));
 NAND4_X2 _31498_ (.A1(_07786_),
    .A2(_07802_),
    .A3(_07818_),
    .A4(_07865_),
    .ZN(_07879_));
 AOI21_X1 _31499_ (.A(_07830_),
    .B1(_07879_),
    .B2(_07781_),
    .ZN(_07880_));
 MUX2_X1 _31500_ (.A(_07880_),
    .B(_07830_),
    .S(_07821_),
    .Z(_07881_));
 AOI21_X1 _31501_ (.A(_07830_),
    .B1(_07879_),
    .B2(_07821_),
    .ZN(_07882_));
 NAND2_X1 _31502_ (.A1(_07781_),
    .A2(_07882_),
    .ZN(_07883_));
 NOR2_X1 _31503_ (.A1(_07830_),
    .A2(_07879_),
    .ZN(_07884_));
 OAI21_X1 _31504_ (.A(_07883_),
    .B1(_07884_),
    .B2(_07781_),
    .ZN(_07885_));
 MUX2_X1 _31505_ (.A(_07881_),
    .B(_07885_),
    .S(_07759_),
    .Z(_07886_));
 NOR2_X1 _31506_ (.A1(_07850_),
    .A2(_07886_),
    .ZN(_00270_));
 CLKBUF_X2 _31507_ (.A(_19749_),
    .Z(_07887_));
 AOI21_X1 _31508_ (.A(_19748_),
    .B1(_07887_),
    .B2(_19750_),
    .ZN(_07888_));
 BUF_X1 _31509_ (.A(_19751_),
    .Z(_07889_));
 NAND2_X1 _31510_ (.A1(_07887_),
    .A2(_07889_),
    .ZN(_07890_));
 CLKBUF_X2 _31511_ (.A(_19754_),
    .Z(_07891_));
 AOI21_X1 _31512_ (.A(_19752_),
    .B1(_19753_),
    .B2(_07891_),
    .ZN(_07892_));
 OAI21_X1 _31513_ (.A(_07888_),
    .B1(_07890_),
    .B2(_07892_),
    .ZN(_07893_));
 INV_X1 _31514_ (.A(_19756_),
    .ZN(_07894_));
 BUF_X1 _31515_ (.A(_19758_),
    .Z(_07895_));
 INV_X1 _31516_ (.A(_19760_),
    .ZN(_07896_));
 AOI21_X1 _31517_ (.A(_19762_),
    .B1(_19763_),
    .B2(_19764_),
    .ZN(_07897_));
 INV_X1 _31518_ (.A(_19761_),
    .ZN(_07898_));
 OAI21_X1 _31519_ (.A(_07896_),
    .B1(_07897_),
    .B2(_07898_),
    .ZN(_07899_));
 BUF_X1 _31520_ (.A(_19759_),
    .Z(_07900_));
 AOI21_X1 _31521_ (.A(_07895_),
    .B1(_07899_),
    .B2(_07900_),
    .ZN(_07901_));
 INV_X1 _31522_ (.A(_19757_),
    .ZN(_07902_));
 OAI21_X2 _31523_ (.A(_07894_),
    .B1(_07901_),
    .B2(_07902_),
    .ZN(_07903_));
 INV_X1 _31524_ (.A(_19753_),
    .ZN(_07904_));
 CLKBUF_X2 _31525_ (.A(_19755_),
    .Z(_07905_));
 INV_X1 _31526_ (.A(_07905_),
    .ZN(_07906_));
 NOR3_X2 _31527_ (.A1(_07904_),
    .A2(_07906_),
    .A3(_07890_),
    .ZN(_07907_));
 AOI21_X2 _31528_ (.A(_07893_),
    .B1(_07903_),
    .B2(_07907_),
    .ZN(_07908_));
 XNOR2_X2 _31529_ (.A(_19747_),
    .B(_07908_),
    .ZN(_07909_));
 INV_X1 _31530_ (.A(_07909_),
    .ZN(_07910_));
 INV_X1 _31531_ (.A(_19752_),
    .ZN(_07911_));
 AOI21_X1 _31532_ (.A(_07891_),
    .B1(_07905_),
    .B2(_07903_),
    .ZN(_07912_));
 OAI21_X2 _31533_ (.A(_07911_),
    .B1(_07912_),
    .B2(_07904_),
    .ZN(_07913_));
 XNOR2_X1 _31534_ (.A(_07889_),
    .B(_07913_),
    .ZN(_07914_));
 XNOR2_X1 _31535_ (.A(_07906_),
    .B(_07903_),
    .ZN(_07915_));
 INV_X1 _31536_ (.A(_19746_),
    .ZN(_07916_));
 INV_X1 _31537_ (.A(_19747_),
    .ZN(_07917_));
 AOI21_X1 _31538_ (.A(_19750_),
    .B1(_07889_),
    .B2(_19752_),
    .ZN(_07918_));
 INV_X1 _31539_ (.A(_07918_),
    .ZN(_07919_));
 AOI21_X1 _31540_ (.A(_19748_),
    .B1(_07919_),
    .B2(_07887_),
    .ZN(_07920_));
 OAI21_X1 _31541_ (.A(_07916_),
    .B1(_07917_),
    .B2(_07920_),
    .ZN(_07921_));
 INV_X1 _31542_ (.A(_07887_),
    .ZN(_07922_));
 NAND2_X1 _31543_ (.A1(_07889_),
    .A2(_19753_),
    .ZN(_07923_));
 NOR3_X2 _31544_ (.A1(_07917_),
    .A2(_07922_),
    .A3(_07923_),
    .ZN(_07924_));
 AOI21_X2 _31545_ (.A(_07891_),
    .B1(_07905_),
    .B2(_19756_),
    .ZN(_07925_));
 OAI21_X1 _31546_ (.A(_07896_),
    .B1(_07898_),
    .B2(_14307_),
    .ZN(_07926_));
 AOI21_X1 _31547_ (.A(_07895_),
    .B1(_07926_),
    .B2(_07900_),
    .ZN(_07927_));
 NAND2_X1 _31548_ (.A1(_07905_),
    .A2(_19757_),
    .ZN(_07928_));
 NOR2_X1 _31549_ (.A1(_07927_),
    .A2(_07928_),
    .ZN(_07929_));
 INV_X1 _31550_ (.A(_07929_),
    .ZN(_07930_));
 NAND2_X1 _31551_ (.A1(_07925_),
    .A2(_07930_),
    .ZN(_07931_));
 AOI21_X1 _31552_ (.A(_07921_),
    .B1(_07924_),
    .B2(_07931_),
    .ZN(_07932_));
 XNOR2_X1 _31553_ (.A(_19745_),
    .B(_07932_),
    .ZN(_19780_));
 AOI21_X1 _31554_ (.A(_07906_),
    .B1(_07902_),
    .B2(_07894_),
    .ZN(_07933_));
 NOR2_X1 _31555_ (.A1(_07891_),
    .A2(_07933_),
    .ZN(_07934_));
 XNOR2_X1 _31556_ (.A(_07904_),
    .B(_07934_),
    .ZN(_07935_));
 XNOR2_X1 _31557_ (.A(_14307_),
    .B(_19761_),
    .ZN(_07936_));
 NOR4_X1 _31558_ (.A1(_14308_),
    .A2(\g_row[1].g_col[1].mult.adder.a[0] ),
    .A3(_19765_),
    .A4(_07936_),
    .ZN(_07937_));
 XNOR2_X1 _31559_ (.A(_07902_),
    .B(_07927_),
    .ZN(_07938_));
 XNOR2_X1 _31560_ (.A(_07900_),
    .B(_07899_),
    .ZN(_07939_));
 NAND4_X1 _31561_ (.A1(_07935_),
    .A2(_07937_),
    .A3(_07938_),
    .A4(_07939_),
    .ZN(_07940_));
 OAI21_X1 _31562_ (.A(_07918_),
    .B1(_07923_),
    .B2(_07925_),
    .ZN(_07941_));
 NOR2_X1 _31563_ (.A1(_07923_),
    .A2(_07930_),
    .ZN(_07942_));
 NOR2_X1 _31564_ (.A1(_07941_),
    .A2(_07942_),
    .ZN(_07943_));
 XNOR2_X1 _31565_ (.A(_07887_),
    .B(_07943_),
    .ZN(_07944_));
 NOR4_X1 _31566_ (.A1(_07915_),
    .A2(_19780_),
    .A3(_07940_),
    .A4(_07944_),
    .ZN(_07945_));
 AND2_X1 _31567_ (.A1(_07914_),
    .A2(_07945_),
    .ZN(_07946_));
 NOR2_X1 _31568_ (.A1(_07910_),
    .A2(_07946_),
    .ZN(_19779_));
 INV_X1 _31569_ (.A(_19726_),
    .ZN(_07947_));
 INV_X1 _31570_ (.A(_19727_),
    .ZN(_07948_));
 INV_X1 _31571_ (.A(_19730_),
    .ZN(_07949_));
 INV_X1 _31572_ (.A(_19731_),
    .ZN(_07950_));
 INV_X1 _31573_ (.A(_19736_),
    .ZN(_07951_));
 BUF_X2 _31574_ (.A(_19739_),
    .Z(_07952_));
 AOI21_X2 _31575_ (.A(_19738_),
    .B1(_07952_),
    .B2(_19740_),
    .ZN(_07953_));
 CLKBUF_X2 _31576_ (.A(_19737_),
    .Z(_07954_));
 INV_X1 _31577_ (.A(_07954_),
    .ZN(_07955_));
 OAI21_X1 _31578_ (.A(_07951_),
    .B1(_07953_),
    .B2(_07955_),
    .ZN(_07956_));
 AOI21_X1 _31579_ (.A(_19734_),
    .B1(_19735_),
    .B2(_07956_),
    .ZN(_07957_));
 BUF_X2 _31580_ (.A(_19743_),
    .Z(_07958_));
 AND2_X1 _31581_ (.A1(_07958_),
    .A2(_19745_),
    .ZN(_07959_));
 AOI21_X1 _31582_ (.A(_19748_),
    .B1(_07941_),
    .B2(_07887_),
    .ZN(_07960_));
 OAI21_X1 _31583_ (.A(_07916_),
    .B1(_07917_),
    .B2(_07960_),
    .ZN(_07961_));
 AOI221_X2 _31584_ (.A(_19742_),
    .B1(_07958_),
    .B2(_19744_),
    .C1(_07959_),
    .C2(_07961_),
    .ZN(_07962_));
 BUF_X2 _31585_ (.A(_19741_),
    .Z(_07963_));
 NAND4_X1 _31586_ (.A1(_19735_),
    .A2(_07954_),
    .A3(_07952_),
    .A4(_07963_),
    .ZN(_07964_));
 OAI21_X1 _31587_ (.A(_07957_),
    .B1(_07962_),
    .B2(_07964_),
    .ZN(_07965_));
 BUF_X2 _31588_ (.A(_19733_),
    .Z(_07966_));
 AOI21_X1 _31589_ (.A(_19732_),
    .B1(_07965_),
    .B2(_07966_),
    .ZN(_07967_));
 OAI21_X1 _31590_ (.A(_07949_),
    .B1(_07950_),
    .B2(_07967_),
    .ZN(_07968_));
 AOI21_X1 _31591_ (.A(_19728_),
    .B1(_19729_),
    .B2(_07968_),
    .ZN(_07969_));
 OAI21_X2 _31592_ (.A(_07947_),
    .B1(_07948_),
    .B2(_07969_),
    .ZN(_07970_));
 INV_X1 _31593_ (.A(_19738_),
    .ZN(_07971_));
 INV_X1 _31594_ (.A(_07952_),
    .ZN(_07972_));
 AOI21_X1 _31595_ (.A(_19740_),
    .B1(_07963_),
    .B2(_19742_),
    .ZN(_07973_));
 OAI21_X1 _31596_ (.A(_07971_),
    .B1(_07972_),
    .B2(_07973_),
    .ZN(_07974_));
 AOI21_X1 _31597_ (.A(_19736_),
    .B1(_07974_),
    .B2(_07954_),
    .ZN(_07975_));
 NAND4_X1 _31598_ (.A1(_07954_),
    .A2(_07952_),
    .A3(_07963_),
    .A4(_07958_),
    .ZN(_07976_));
 AOI21_X1 _31599_ (.A(_19744_),
    .B1(_19745_),
    .B2(_19746_),
    .ZN(_07977_));
 NAND2_X1 _31600_ (.A1(_19745_),
    .A2(_19747_),
    .ZN(_07978_));
 OAI21_X1 _31601_ (.A(_07977_),
    .B1(_07978_),
    .B2(_07888_),
    .ZN(_07979_));
 NOR2_X1 _31602_ (.A1(_07890_),
    .A2(_07978_),
    .ZN(_07980_));
 INV_X1 _31603_ (.A(_07895_),
    .ZN(_07981_));
 OAI21_X1 _31604_ (.A(_07894_),
    .B1(_07981_),
    .B2(_07902_),
    .ZN(_07982_));
 AOI21_X1 _31605_ (.A(_07891_),
    .B1(_07905_),
    .B2(_07982_),
    .ZN(_07983_));
 OAI21_X1 _31606_ (.A(_07911_),
    .B1(_07983_),
    .B2(_07904_),
    .ZN(_07984_));
 AOI21_X1 _31607_ (.A(_07979_),
    .B1(_07980_),
    .B2(_07984_),
    .ZN(_07985_));
 OAI21_X1 _31608_ (.A(_07975_),
    .B1(_07976_),
    .B2(_07985_),
    .ZN(_07986_));
 AOI21_X1 _31609_ (.A(_19734_),
    .B1(_19735_),
    .B2(_07986_),
    .ZN(_07987_));
 INV_X1 _31610_ (.A(_07987_),
    .ZN(_07988_));
 AOI21_X1 _31611_ (.A(_19732_),
    .B1(_07988_),
    .B2(_07966_),
    .ZN(_07989_));
 OAI21_X1 _31612_ (.A(_07949_),
    .B1(_07950_),
    .B2(_07989_),
    .ZN(_07990_));
 AOI21_X2 _31613_ (.A(_19728_),
    .B1(_19729_),
    .B2(_07990_),
    .ZN(_07991_));
 XNOR2_X2 _31614_ (.A(_19727_),
    .B(_07991_),
    .ZN(_07992_));
 NAND2_X1 _31615_ (.A1(_07924_),
    .A2(_07959_),
    .ZN(_07993_));
 OAI21_X2 _31616_ (.A(_07962_),
    .B1(_07993_),
    .B2(_07930_),
    .ZN(_07994_));
 INV_X1 _31617_ (.A(_07994_),
    .ZN(_07995_));
 OAI21_X1 _31618_ (.A(_07957_),
    .B1(_07964_),
    .B2(_07995_),
    .ZN(_07996_));
 XOR2_X2 _31619_ (.A(_07966_),
    .B(_07996_),
    .Z(_07997_));
 INV_X1 _31620_ (.A(_19734_),
    .ZN(_07998_));
 INV_X1 _31621_ (.A(_19735_),
    .ZN(_07999_));
 NAND2_X1 _31622_ (.A1(_07963_),
    .A2(_07958_),
    .ZN(_08000_));
 OAI21_X1 _31623_ (.A(_07973_),
    .B1(_08000_),
    .B2(_07977_),
    .ZN(_08001_));
 INV_X1 _31624_ (.A(_19762_),
    .ZN(_08002_));
 OAI21_X1 _31625_ (.A(_07896_),
    .B1(_08002_),
    .B2(_07898_),
    .ZN(_08003_));
 AOI21_X1 _31626_ (.A(_07895_),
    .B1(_08003_),
    .B2(_07900_),
    .ZN(_08004_));
 OAI21_X1 _31627_ (.A(_07894_),
    .B1(_08004_),
    .B2(_07902_),
    .ZN(_08005_));
 AOI21_X1 _31628_ (.A(_07893_),
    .B1(_07907_),
    .B2(_08005_),
    .ZN(_08006_));
 NOR3_X1 _31629_ (.A1(_08000_),
    .A2(_07978_),
    .A3(_08006_),
    .ZN(_08007_));
 OAI21_X1 _31630_ (.A(_07952_),
    .B1(_08001_),
    .B2(_08007_),
    .ZN(_08008_));
 NAND2_X1 _31631_ (.A1(_07971_),
    .A2(_08008_),
    .ZN(_08009_));
 AOI21_X1 _31632_ (.A(_19736_),
    .B1(_08009_),
    .B2(_07954_),
    .ZN(_08010_));
 OAI21_X1 _31633_ (.A(_07998_),
    .B1(_07999_),
    .B2(_08010_),
    .ZN(_08011_));
 AOI21_X2 _31634_ (.A(_19732_),
    .B1(_08011_),
    .B2(_07966_),
    .ZN(_08012_));
 XNOR2_X2 _31635_ (.A(_19731_),
    .B(_08012_),
    .ZN(_08013_));
 AOI21_X2 _31636_ (.A(_19742_),
    .B1(_07958_),
    .B2(_19744_),
    .ZN(_08014_));
 NAND2_X1 _31637_ (.A1(_07952_),
    .A2(_07963_),
    .ZN(_08015_));
 NAND3_X1 _31638_ (.A1(_07952_),
    .A2(_07963_),
    .A3(_07959_),
    .ZN(_08016_));
 OAI221_X2 _31639_ (.A(_07953_),
    .B1(_08014_),
    .B2(_08015_),
    .C1(_08016_),
    .C2(_07932_),
    .ZN(_08017_));
 XNOR2_X2 _31640_ (.A(_07955_),
    .B(_08017_),
    .ZN(_08018_));
 AOI21_X2 _31641_ (.A(_07979_),
    .B1(_07980_),
    .B2(_07913_),
    .ZN(_08019_));
 XNOR2_X2 _31642_ (.A(_07958_),
    .B(_08019_),
    .ZN(_08020_));
 AND3_X1 _31643_ (.A1(_07909_),
    .A2(_19780_),
    .A3(_08020_),
    .ZN(_08021_));
 NOR3_X1 _31644_ (.A1(_07908_),
    .A2(_08000_),
    .A3(_07978_),
    .ZN(_08022_));
 NOR2_X1 _31645_ (.A1(_08001_),
    .A2(_08022_),
    .ZN(_08023_));
 XNOR2_X2 _31646_ (.A(_07972_),
    .B(_08023_),
    .ZN(_08024_));
 INV_X1 _31647_ (.A(_08024_),
    .ZN(_08025_));
 XOR2_X2 _31648_ (.A(_07963_),
    .B(_07994_),
    .Z(_08026_));
 AND3_X1 _31649_ (.A1(_08021_),
    .A2(_08025_),
    .A3(_08026_),
    .ZN(_08027_));
 OAI21_X1 _31650_ (.A(_07975_),
    .B1(_07976_),
    .B2(_08019_),
    .ZN(_08028_));
 XNOR2_X2 _31651_ (.A(_07999_),
    .B(_08028_),
    .ZN(_08029_));
 NAND3_X1 _31652_ (.A1(_08018_),
    .A2(_08027_),
    .A3(_08029_),
    .ZN(_08030_));
 INV_X1 _31653_ (.A(_08030_),
    .ZN(_08031_));
 NAND3_X1 _31654_ (.A1(_07997_),
    .A2(_08013_),
    .A3(_08031_),
    .ZN(_08032_));
 AOI21_X1 _31655_ (.A(_07895_),
    .B1(_19760_),
    .B2(_07900_),
    .ZN(_08033_));
 OAI21_X1 _31656_ (.A(_07925_),
    .B1(_07928_),
    .B2(_08033_),
    .ZN(_08034_));
 AOI21_X1 _31657_ (.A(_07921_),
    .B1(_07924_),
    .B2(_08034_),
    .ZN(_08035_));
 OAI221_X1 _31658_ (.A(_07953_),
    .B1(_08014_),
    .B2(_08015_),
    .C1(_08016_),
    .C2(_08035_),
    .ZN(_08036_));
 AOI21_X1 _31659_ (.A(_19736_),
    .B1(_08036_),
    .B2(_07954_),
    .ZN(_08037_));
 OAI21_X1 _31660_ (.A(_07998_),
    .B1(_07999_),
    .B2(_08037_),
    .ZN(_08038_));
 AOI21_X1 _31661_ (.A(_19732_),
    .B1(_08038_),
    .B2(_07966_),
    .ZN(_08039_));
 OAI21_X1 _31662_ (.A(_07949_),
    .B1(_07950_),
    .B2(_08039_),
    .ZN(_08040_));
 XNOR2_X2 _31663_ (.A(_19729_),
    .B(_08040_),
    .ZN(_08041_));
 OR2_X1 _31664_ (.A1(_08032_),
    .A2(_08041_),
    .ZN(_08042_));
 INV_X1 _31665_ (.A(_08042_),
    .ZN(_08043_));
 NAND2_X1 _31666_ (.A1(_07992_),
    .A2(_08043_),
    .ZN(_08044_));
 XNOR2_X1 _31667_ (.A(_07970_),
    .B(_08044_),
    .ZN(_08045_));
 BUF_X1 _31668_ (.A(_08045_),
    .Z(_14310_));
 INV_X1 _31669_ (.A(_14310_),
    .ZN(_14314_));
 OR4_X1 _31670_ (.A1(\g_row[1].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08046_));
 OAI21_X2 _31671_ (.A(_07176_),
    .B1(_08046_),
    .B2(\g_row[1].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08047_));
 AND4_X1 _31672_ (.A1(\g_row[1].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08048_));
 AOI21_X4 _31673_ (.A(_07180_),
    .B1(_08048_),
    .B2(\g_row[1].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08049_));
 INV_X1 _31674_ (.A(_14312_),
    .ZN(_08050_));
 AOI21_X1 _31675_ (.A(_08047_),
    .B1(_08049_),
    .B2(_08050_),
    .ZN(_00273_));
 INV_X1 _31676_ (.A(_19769_),
    .ZN(_08051_));
 AOI21_X1 _31677_ (.A(_08047_),
    .B1(_08049_),
    .B2(_08051_),
    .ZN(_00274_));
 INV_X1 _31678_ (.A(_14320_),
    .ZN(_08052_));
 AOI21_X1 _31679_ (.A(_08047_),
    .B1(_08049_),
    .B2(_08052_),
    .ZN(_00275_));
 XOR2_X1 _31680_ (.A(_14319_),
    .B(_19778_),
    .Z(_08053_));
 AOI21_X1 _31681_ (.A(_08047_),
    .B1(_08049_),
    .B2(_08053_),
    .ZN(_00276_));
 AOI21_X1 _31682_ (.A(_19773_),
    .B1(_19774_),
    .B2(_19768_),
    .ZN(_08054_));
 INV_X1 _31683_ (.A(_08054_),
    .ZN(_08055_));
 AOI21_X1 _31684_ (.A(_19777_),
    .B1(_08055_),
    .B2(_19778_),
    .ZN(_08056_));
 XNOR2_X1 _31685_ (.A(\g_row[1].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_19775_),
    .ZN(_08057_));
 XNOR2_X1 _31686_ (.A(_07174_),
    .B(_08057_),
    .ZN(_08058_));
 XNOR2_X1 _31687_ (.A(_08056_),
    .B(_08058_),
    .ZN(_08059_));
 AOI21_X1 _31688_ (.A(_08047_),
    .B1(_08049_),
    .B2(_08059_),
    .ZN(_00277_));
 INV_X1 _31689_ (.A(_08047_),
    .ZN(_08060_));
 NAND2_X4 _31690_ (.A1(_08060_),
    .A2(_08049_),
    .ZN(_08061_));
 NAND2_X1 _31691_ (.A1(_19782_),
    .A2(_14310_),
    .ZN(_08062_));
 NAND3_X1 _31692_ (.A1(_07909_),
    .A2(_07946_),
    .A3(_14314_),
    .ZN(_08063_));
 AOI21_X1 _31693_ (.A(_08061_),
    .B1(_08062_),
    .B2(_08063_),
    .ZN(_00272_));
 INV_X1 _31694_ (.A(_19782_),
    .ZN(_08064_));
 XNOR2_X1 _31695_ (.A(_19781_),
    .B(_08020_),
    .ZN(_08065_));
 MUX2_X1 _31696_ (.A(_08064_),
    .B(_08065_),
    .S(_14310_),
    .Z(_08066_));
 NOR2_X1 _31697_ (.A1(_08061_),
    .A2(_08066_),
    .ZN(_00278_));
 XNOR2_X1 _31698_ (.A(_08021_),
    .B(_08026_),
    .ZN(_08067_));
 MUX2_X1 _31699_ (.A(_08065_),
    .B(_08067_),
    .S(_14310_),
    .Z(_08068_));
 NOR2_X1 _31700_ (.A1(_08061_),
    .A2(_08068_),
    .ZN(_00279_));
 NAND3_X1 _31701_ (.A1(_19781_),
    .A2(_08020_),
    .A3(_08026_),
    .ZN(_08069_));
 XNOR2_X1 _31702_ (.A(_08024_),
    .B(_08069_),
    .ZN(_08070_));
 MUX2_X1 _31703_ (.A(_08067_),
    .B(_08070_),
    .S(_14310_),
    .Z(_08071_));
 NOR2_X1 _31704_ (.A1(_08061_),
    .A2(_08071_),
    .ZN(_00280_));
 XNOR2_X1 _31705_ (.A(_08018_),
    .B(_08027_),
    .ZN(_08072_));
 MUX2_X1 _31706_ (.A(_08070_),
    .B(_08072_),
    .S(_14310_),
    .Z(_08073_));
 NOR2_X1 _31707_ (.A1(_08061_),
    .A2(_08073_),
    .ZN(_00281_));
 INV_X1 _31708_ (.A(_08018_),
    .ZN(_08074_));
 NOR3_X1 _31709_ (.A1(_08074_),
    .A2(_08024_),
    .A3(_08069_),
    .ZN(_08075_));
 XNOR2_X1 _31710_ (.A(_08029_),
    .B(_08075_),
    .ZN(_08076_));
 MUX2_X1 _31711_ (.A(_08072_),
    .B(_08076_),
    .S(_14310_),
    .Z(_08077_));
 NOR2_X1 _31712_ (.A1(_08061_),
    .A2(_08077_),
    .ZN(_00282_));
 XOR2_X1 _31713_ (.A(_07997_),
    .B(_08030_),
    .Z(_08078_));
 MUX2_X1 _31714_ (.A(_08076_),
    .B(_08078_),
    .S(_08045_),
    .Z(_08079_));
 NOR2_X1 _31715_ (.A1(_08061_),
    .A2(_08079_),
    .ZN(_00283_));
 NOR2_X1 _31716_ (.A1(_14310_),
    .A2(_08078_),
    .ZN(_08080_));
 NAND3_X1 _31717_ (.A1(_07997_),
    .A2(_08029_),
    .A3(_08075_),
    .ZN(_08081_));
 XNOR2_X1 _31718_ (.A(_08013_),
    .B(_08081_),
    .ZN(_08082_));
 AOI21_X1 _31719_ (.A(_08080_),
    .B1(_08082_),
    .B2(_14310_),
    .ZN(_08083_));
 NOR2_X1 _31720_ (.A1(_08061_),
    .A2(_08083_),
    .ZN(_00284_));
 NOR2_X1 _31721_ (.A1(_08042_),
    .A2(_08082_),
    .ZN(_08084_));
 NAND2_X1 _31722_ (.A1(_08044_),
    .A2(_08082_),
    .ZN(_08085_));
 NAND2_X1 _31723_ (.A1(_08032_),
    .A2(_08041_),
    .ZN(_08086_));
 OAI21_X1 _31724_ (.A(_08086_),
    .B1(_08042_),
    .B2(_07992_),
    .ZN(_08087_));
 MUX2_X1 _31725_ (.A(_08085_),
    .B(_08087_),
    .S(_07970_),
    .Z(_08088_));
 NOR3_X1 _31726_ (.A1(_08061_),
    .A2(_08084_),
    .A3(_08088_),
    .ZN(_00285_));
 NAND4_X2 _31727_ (.A1(_07997_),
    .A2(_08013_),
    .A3(_08029_),
    .A4(_08075_),
    .ZN(_08089_));
 AOI21_X1 _31728_ (.A(_08041_),
    .B1(_08089_),
    .B2(_07992_),
    .ZN(_08090_));
 MUX2_X1 _31729_ (.A(_08090_),
    .B(_08041_),
    .S(_08032_),
    .Z(_08091_));
 AOI21_X1 _31730_ (.A(_08041_),
    .B1(_08089_),
    .B2(_08032_),
    .ZN(_08092_));
 NAND2_X1 _31731_ (.A1(_07992_),
    .A2(_08092_),
    .ZN(_08093_));
 NOR2_X1 _31732_ (.A1(_08041_),
    .A2(_08089_),
    .ZN(_08094_));
 OAI21_X1 _31733_ (.A(_08093_),
    .B1(_08094_),
    .B2(_07992_),
    .ZN(_08095_));
 MUX2_X1 _31734_ (.A(_08091_),
    .B(_08095_),
    .S(_07970_),
    .Z(_08096_));
 NOR2_X1 _31735_ (.A1(_08061_),
    .A2(_08096_),
    .ZN(_00286_));
 BUF_X2 _31736_ (.A(_19804_),
    .Z(_08097_));
 INV_X1 _31737_ (.A(_19805_),
    .ZN(_08098_));
 CLKBUF_X2 _31738_ (.A(_19808_),
    .Z(_08099_));
 INV_X1 _31739_ (.A(_19809_),
    .ZN(_08100_));
 CLKBUF_X2 _31740_ (.A(_19812_),
    .Z(_08101_));
 INV_X1 _31741_ (.A(_19813_),
    .ZN(_08102_));
 BUF_X1 _31742_ (.A(_19815_),
    .Z(_08103_));
 INV_X1 _31743_ (.A(_19817_),
    .ZN(_08104_));
 AOI21_X1 _31744_ (.A(_19819_),
    .B1(_19820_),
    .B2(_19821_),
    .ZN(_08105_));
 INV_X1 _31745_ (.A(_19818_),
    .ZN(_08106_));
 OAI21_X1 _31746_ (.A(_08104_),
    .B1(_08105_),
    .B2(_08106_),
    .ZN(_08107_));
 AOI21_X1 _31747_ (.A(_08103_),
    .B1(_08107_),
    .B2(_19816_),
    .ZN(_08108_));
 BUF_X1 _31748_ (.A(_19814_),
    .Z(_08109_));
 INV_X1 _31749_ (.A(_08109_),
    .ZN(_08110_));
 OAI21_X1 _31750_ (.A(_08102_),
    .B1(_08108_),
    .B2(_08110_),
    .ZN(_08111_));
 AOI21_X1 _31751_ (.A(_19811_),
    .B1(_08101_),
    .B2(_08111_),
    .ZN(_08112_));
 CLKBUF_X2 _31752_ (.A(_19810_),
    .Z(_08113_));
 INV_X1 _31753_ (.A(_08113_),
    .ZN(_08114_));
 OAI21_X1 _31754_ (.A(_08100_),
    .B1(_08112_),
    .B2(_08114_),
    .ZN(_08115_));
 AOI21_X1 _31755_ (.A(_19807_),
    .B1(_08099_),
    .B2(_08115_),
    .ZN(_08116_));
 BUF_X2 _31756_ (.A(_19806_),
    .Z(_08117_));
 INV_X1 _31757_ (.A(_08117_),
    .ZN(_08118_));
 OAI21_X1 _31758_ (.A(_08098_),
    .B1(_08116_),
    .B2(_08118_),
    .ZN(_08119_));
 XNOR2_X1 _31759_ (.A(_08097_),
    .B(_08119_),
    .ZN(_08120_));
 INV_X1 _31760_ (.A(_08099_),
    .ZN(_08121_));
 XNOR2_X1 _31761_ (.A(_08121_),
    .B(_08115_),
    .ZN(_08122_));
 BUF_X1 _31762_ (.A(_19802_),
    .Z(_08123_));
 INV_X1 _31763_ (.A(_08123_),
    .ZN(_08124_));
 AOI21_X1 _31764_ (.A(_19807_),
    .B1(_08099_),
    .B2(_19809_),
    .ZN(_08125_));
 OAI21_X1 _31765_ (.A(_08098_),
    .B1(_08125_),
    .B2(_08118_),
    .ZN(_08126_));
 AOI21_X1 _31766_ (.A(_19803_),
    .B1(_08097_),
    .B2(_08126_),
    .ZN(_08127_));
 NAND4_X2 _31767_ (.A1(_08097_),
    .A2(_08117_),
    .A3(_08099_),
    .A4(_08113_),
    .ZN(_08128_));
 AOI21_X2 _31768_ (.A(_19811_),
    .B1(_08101_),
    .B2(_19813_),
    .ZN(_08129_));
 OAI21_X1 _31769_ (.A(_08104_),
    .B1(_08106_),
    .B2(_14324_),
    .ZN(_08130_));
 AOI21_X1 _31770_ (.A(_08103_),
    .B1(_08130_),
    .B2(_19816_),
    .ZN(_08131_));
 NAND2_X1 _31771_ (.A1(_08101_),
    .A2(_08109_),
    .ZN(_08132_));
 OR2_X1 _31772_ (.A1(_08131_),
    .A2(_08132_),
    .ZN(_08133_));
 AND2_X1 _31773_ (.A1(_08129_),
    .A2(_08133_),
    .ZN(_08134_));
 OAI21_X2 _31774_ (.A(_08127_),
    .B1(_08128_),
    .B2(_08134_),
    .ZN(_08135_));
 XNOR2_X2 _31775_ (.A(_08124_),
    .B(_08135_),
    .ZN(_19836_));
 XNOR2_X1 _31776_ (.A(_08101_),
    .B(_08111_),
    .ZN(_08136_));
 NAND2_X1 _31777_ (.A1(_08099_),
    .A2(_08113_),
    .ZN(_08137_));
 OAI21_X1 _31778_ (.A(_08125_),
    .B1(_08137_),
    .B2(_08129_),
    .ZN(_08138_));
 INV_X1 _31779_ (.A(_08138_),
    .ZN(_08139_));
 OAI21_X1 _31780_ (.A(_08139_),
    .B1(_08133_),
    .B2(_08137_),
    .ZN(_08140_));
 XNOR2_X1 _31781_ (.A(_08117_),
    .B(_08140_),
    .ZN(_08141_));
 XNOR2_X1 _31782_ (.A(_14324_),
    .B(_19818_),
    .ZN(_08142_));
 OR4_X1 _31783_ (.A1(_14325_),
    .A2(\g_row[1].g_col[2].mult.adder.a[0] ),
    .A3(_19822_),
    .A4(_08142_),
    .ZN(_08143_));
 XNOR2_X1 _31784_ (.A(_08109_),
    .B(_08131_),
    .ZN(_08144_));
 INV_X1 _31785_ (.A(_19816_),
    .ZN(_08145_));
 XNOR2_X1 _31786_ (.A(_08145_),
    .B(_08107_),
    .ZN(_08146_));
 NOR3_X1 _31787_ (.A1(_08143_),
    .A2(_08144_),
    .A3(_08146_),
    .ZN(_08147_));
 XNOR2_X1 _31788_ (.A(_08114_),
    .B(_08134_),
    .ZN(_08148_));
 NAND4_X1 _31789_ (.A1(_08136_),
    .A2(_08141_),
    .A3(_08147_),
    .A4(_08148_),
    .ZN(_08149_));
 NOR3_X1 _31790_ (.A1(_08122_),
    .A2(_19836_),
    .A3(_08149_),
    .ZN(_08150_));
 NOR2_X1 _31791_ (.A1(_08120_),
    .A2(_08150_),
    .ZN(_19837_));
 INV_X1 _31792_ (.A(_19783_),
    .ZN(_08151_));
 INV_X1 _31793_ (.A(_19784_),
    .ZN(_08152_));
 INV_X1 _31794_ (.A(_19787_),
    .ZN(_08153_));
 INV_X1 _31795_ (.A(_19788_),
    .ZN(_08154_));
 BUF_X2 _31796_ (.A(_19792_),
    .Z(_08155_));
 INV_X1 _31797_ (.A(_19793_),
    .ZN(_08156_));
 CLKBUF_X2 _31798_ (.A(_19796_),
    .Z(_08157_));
 AOI21_X1 _31799_ (.A(_19795_),
    .B1(_08157_),
    .B2(_19797_),
    .ZN(_08158_));
 CLKBUF_X3 _31800_ (.A(_19794_),
    .Z(_08159_));
 INV_X1 _31801_ (.A(_08159_),
    .ZN(_08160_));
 OAI21_X1 _31802_ (.A(_08156_),
    .B1(_08158_),
    .B2(_08160_),
    .ZN(_08161_));
 AOI21_X1 _31803_ (.A(_19791_),
    .B1(_08155_),
    .B2(_08161_),
    .ZN(_08162_));
 BUF_X2 _31804_ (.A(_19800_),
    .Z(_08163_));
 AOI21_X1 _31805_ (.A(_19799_),
    .B1(_08163_),
    .B2(_19801_),
    .ZN(_08164_));
 INV_X1 _31806_ (.A(_19803_),
    .ZN(_08165_));
 INV_X1 _31807_ (.A(_08097_),
    .ZN(_08166_));
 AOI21_X1 _31808_ (.A(_19805_),
    .B1(_08138_),
    .B2(_08117_),
    .ZN(_08167_));
 OAI21_X1 _31809_ (.A(_08165_),
    .B1(_08166_),
    .B2(_08167_),
    .ZN(_08168_));
 NAND3_X1 _31810_ (.A1(_08163_),
    .A2(_08123_),
    .A3(_08168_),
    .ZN(_08169_));
 AND2_X1 _31811_ (.A1(_08164_),
    .A2(_08169_),
    .ZN(_08170_));
 BUF_X2 _31812_ (.A(_19798_),
    .Z(_08171_));
 AND2_X1 _31813_ (.A1(_08157_),
    .A2(_08171_),
    .ZN(_08172_));
 NAND3_X1 _31814_ (.A1(_08155_),
    .A2(_08159_),
    .A3(_08172_),
    .ZN(_08173_));
 OAI21_X1 _31815_ (.A(_08162_),
    .B1(_08170_),
    .B2(_08173_),
    .ZN(_08174_));
 CLKBUF_X2 _31816_ (.A(_19790_),
    .Z(_08175_));
 AOI21_X1 _31817_ (.A(_19789_),
    .B1(_08174_),
    .B2(_08175_),
    .ZN(_08176_));
 OAI21_X1 _31818_ (.A(_08153_),
    .B1(_08154_),
    .B2(_08176_),
    .ZN(_08177_));
 AOI21_X2 _31819_ (.A(_19785_),
    .B1(_19786_),
    .B2(_08177_),
    .ZN(_08178_));
 OAI21_X2 _31820_ (.A(_08151_),
    .B1(_08152_),
    .B2(_08178_),
    .ZN(_08179_));
 INV_X1 _31821_ (.A(_19789_),
    .ZN(_08180_));
 AOI21_X2 _31822_ (.A(_19797_),
    .B1(_08171_),
    .B2(_19799_),
    .ZN(_08181_));
 NAND2_X1 _31823_ (.A1(_08171_),
    .A2(_08163_),
    .ZN(_08182_));
 INV_X1 _31824_ (.A(_19807_),
    .ZN(_08183_));
 INV_X1 _31825_ (.A(_19811_),
    .ZN(_08184_));
 INV_X1 _31826_ (.A(_08101_),
    .ZN(_08185_));
 INV_X1 _31827_ (.A(_08103_),
    .ZN(_08186_));
 AOI21_X1 _31828_ (.A(_19817_),
    .B1(_19819_),
    .B2(_19818_),
    .ZN(_08187_));
 OAI21_X1 _31829_ (.A(_08186_),
    .B1(_08187_),
    .B2(_08145_),
    .ZN(_08188_));
 AOI21_X1 _31830_ (.A(_19813_),
    .B1(_08188_),
    .B2(_08109_),
    .ZN(_08189_));
 OAI21_X1 _31831_ (.A(_08184_),
    .B1(_08185_),
    .B2(_08189_),
    .ZN(_08190_));
 AOI21_X1 _31832_ (.A(_19809_),
    .B1(_08190_),
    .B2(_08113_),
    .ZN(_08191_));
 OAI21_X1 _31833_ (.A(_08183_),
    .B1(_08121_),
    .B2(_08191_),
    .ZN(_08192_));
 AOI21_X1 _31834_ (.A(_19805_),
    .B1(_08192_),
    .B2(_08117_),
    .ZN(_08193_));
 OAI21_X1 _31835_ (.A(_08165_),
    .B1(_08166_),
    .B2(_08193_),
    .ZN(_08194_));
 AOI21_X1 _31836_ (.A(_19801_),
    .B1(_08194_),
    .B2(_08123_),
    .ZN(_08195_));
 OAI21_X1 _31837_ (.A(_08181_),
    .B1(_08182_),
    .B2(_08195_),
    .ZN(_08196_));
 AOI21_X1 _31838_ (.A(_19795_),
    .B1(_08157_),
    .B2(_08196_),
    .ZN(_08197_));
 OAI21_X1 _31839_ (.A(_08156_),
    .B1(_08197_),
    .B2(_08160_),
    .ZN(_08198_));
 AOI21_X1 _31840_ (.A(_19791_),
    .B1(_08155_),
    .B2(_08198_),
    .ZN(_08199_));
 INV_X1 _31841_ (.A(_08175_),
    .ZN(_08200_));
 OAI21_X1 _31842_ (.A(_08180_),
    .B1(_08199_),
    .B2(_08200_),
    .ZN(_08201_));
 XNOR2_X2 _31843_ (.A(_19788_),
    .B(_08201_),
    .ZN(_08202_));
 INV_X1 _31844_ (.A(_08157_),
    .ZN(_08203_));
 INV_X1 _31845_ (.A(_19801_),
    .ZN(_08204_));
 AOI21_X1 _31846_ (.A(_19803_),
    .B1(_08097_),
    .B2(_08119_),
    .ZN(_08205_));
 OAI21_X1 _31847_ (.A(_08204_),
    .B1(_08205_),
    .B2(_08124_),
    .ZN(_08206_));
 NAND3_X1 _31848_ (.A1(_08171_),
    .A2(_08163_),
    .A3(_08206_),
    .ZN(_08207_));
 NAND2_X1 _31849_ (.A1(_08181_),
    .A2(_08207_),
    .ZN(_08208_));
 XNOR2_X1 _31850_ (.A(_08203_),
    .B(_08208_),
    .ZN(_08209_));
 XNOR2_X2 _31851_ (.A(_08163_),
    .B(_08206_),
    .ZN(_08210_));
 XNOR2_X1 _31852_ (.A(_08166_),
    .B(_08119_),
    .ZN(_08211_));
 NAND2_X1 _31853_ (.A1(_08211_),
    .A2(_19836_),
    .ZN(_08212_));
 NOR2_X1 _31854_ (.A1(_08210_),
    .A2(_08212_),
    .ZN(_08213_));
 NAND2_X1 _31855_ (.A1(_08163_),
    .A2(_08123_),
    .ZN(_08214_));
 OR2_X1 _31856_ (.A1(_08128_),
    .A2(_08214_),
    .ZN(_08215_));
 OAI21_X2 _31857_ (.A(_08170_),
    .B1(_08215_),
    .B2(_08133_),
    .ZN(_08216_));
 XOR2_X2 _31858_ (.A(_08171_),
    .B(_08216_),
    .Z(_08217_));
 AND3_X1 _31859_ (.A1(_08209_),
    .A2(_08213_),
    .A3(_08217_),
    .ZN(_08218_));
 NAND2_X1 _31860_ (.A1(_08157_),
    .A2(_08171_),
    .ZN(_08219_));
 OAI21_X1 _31861_ (.A(_08158_),
    .B1(_08164_),
    .B2(_08219_),
    .ZN(_08220_));
 NOR2_X1 _31862_ (.A1(_08214_),
    .A2(_08219_),
    .ZN(_08221_));
 AOI21_X2 _31863_ (.A(_08220_),
    .B1(_08221_),
    .B2(_08135_),
    .ZN(_08222_));
 XNOR2_X2 _31864_ (.A(_08159_),
    .B(_08222_),
    .ZN(_08223_));
 NOR3_X1 _31865_ (.A1(_08160_),
    .A2(_08203_),
    .A3(_08182_),
    .ZN(_08224_));
 INV_X1 _31866_ (.A(_19795_),
    .ZN(_08225_));
 OAI21_X1 _31867_ (.A(_08225_),
    .B1(_08203_),
    .B2(_08181_),
    .ZN(_08226_));
 AOI221_X2 _31868_ (.A(_19793_),
    .B1(_08206_),
    .B2(_08224_),
    .C1(_08226_),
    .C2(_08159_),
    .ZN(_08227_));
 XNOR2_X2 _31869_ (.A(_08155_),
    .B(_08227_),
    .ZN(_08228_));
 NAND3_X1 _31870_ (.A1(_08218_),
    .A2(_08223_),
    .A3(_08228_),
    .ZN(_08229_));
 NAND4_X1 _31871_ (.A1(_08155_),
    .A2(_08159_),
    .A3(_08172_),
    .A4(_08216_),
    .ZN(_08230_));
 NAND2_X1 _31872_ (.A1(_08162_),
    .A2(_08230_),
    .ZN(_08231_));
 XNOR2_X2 _31873_ (.A(_08175_),
    .B(_08231_),
    .ZN(_08232_));
 NOR3_X1 _31874_ (.A1(_08202_),
    .A2(_08229_),
    .A3(_08232_),
    .ZN(_08233_));
 INV_X1 _31875_ (.A(_19785_),
    .ZN(_08234_));
 INV_X1 _31876_ (.A(_19786_),
    .ZN(_08235_));
 AOI21_X1 _31877_ (.A(_19793_),
    .B1(_08226_),
    .B2(_08159_),
    .ZN(_08236_));
 NAND4_X1 _31878_ (.A1(_08159_),
    .A2(_08157_),
    .A3(_08171_),
    .A4(_08163_),
    .ZN(_08237_));
 AOI21_X1 _31879_ (.A(_19813_),
    .B1(_08103_),
    .B2(_08109_),
    .ZN(_08238_));
 OAI21_X1 _31880_ (.A(_08184_),
    .B1(_08185_),
    .B2(_08238_),
    .ZN(_08239_));
 AOI21_X1 _31881_ (.A(_19809_),
    .B1(_08239_),
    .B2(_08113_),
    .ZN(_08240_));
 OAI21_X1 _31882_ (.A(_08183_),
    .B1(_08121_),
    .B2(_08240_),
    .ZN(_08241_));
 AOI21_X1 _31883_ (.A(_19805_),
    .B1(_08241_),
    .B2(_08117_),
    .ZN(_08242_));
 OAI21_X1 _31884_ (.A(_08165_),
    .B1(_08166_),
    .B2(_08242_),
    .ZN(_08243_));
 AOI21_X1 _31885_ (.A(_19801_),
    .B1(_08243_),
    .B2(_08123_),
    .ZN(_08244_));
 OAI21_X1 _31886_ (.A(_08236_),
    .B1(_08237_),
    .B2(_08244_),
    .ZN(_08245_));
 AOI21_X1 _31887_ (.A(_19791_),
    .B1(_08155_),
    .B2(_08245_),
    .ZN(_08246_));
 OAI21_X1 _31888_ (.A(_08180_),
    .B1(_08246_),
    .B2(_08200_),
    .ZN(_08247_));
 AOI21_X1 _31889_ (.A(_19787_),
    .B1(_19788_),
    .B2(_08247_),
    .ZN(_08248_));
 OAI21_X1 _31890_ (.A(_08234_),
    .B1(_08235_),
    .B2(_08248_),
    .ZN(_08249_));
 XNOR2_X2 _31891_ (.A(_19784_),
    .B(_08249_),
    .ZN(_08250_));
 INV_X1 _31892_ (.A(_08155_),
    .ZN(_08251_));
 NOR3_X1 _31893_ (.A1(_08166_),
    .A2(_08118_),
    .A3(_08137_),
    .ZN(_08252_));
 AOI21_X1 _31894_ (.A(_08103_),
    .B1(_19817_),
    .B2(_19816_),
    .ZN(_08253_));
 OAI21_X1 _31895_ (.A(_08129_),
    .B1(_08132_),
    .B2(_08253_),
    .ZN(_08254_));
 AOI221_X2 _31896_ (.A(_19803_),
    .B1(_08097_),
    .B2(_08126_),
    .C1(_08252_),
    .C2(_08254_),
    .ZN(_08255_));
 NOR3_X1 _31897_ (.A1(_08214_),
    .A2(_08219_),
    .A3(_08255_),
    .ZN(_08256_));
 OAI21_X1 _31898_ (.A(_08159_),
    .B1(_08220_),
    .B2(_08256_),
    .ZN(_08257_));
 AOI21_X1 _31899_ (.A(_08251_),
    .B1(_08156_),
    .B2(_08257_),
    .ZN(_08258_));
 OAI21_X1 _31900_ (.A(_08175_),
    .B1(_08258_),
    .B2(_19791_),
    .ZN(_08259_));
 AOI21_X1 _31901_ (.A(_08154_),
    .B1(_08180_),
    .B2(_08259_),
    .ZN(_08260_));
 NOR2_X1 _31902_ (.A1(_19787_),
    .A2(_08260_),
    .ZN(_08261_));
 XNOR2_X2 _31903_ (.A(_08235_),
    .B(_08261_),
    .ZN(_08262_));
 NOR2_X1 _31904_ (.A1(_08250_),
    .A2(_08262_),
    .ZN(_08263_));
 NAND2_X1 _31905_ (.A1(_08233_),
    .A2(_08263_),
    .ZN(_08264_));
 XNOR2_X1 _31906_ (.A(_08179_),
    .B(_08264_),
    .ZN(_14327_));
 INV_X1 _31907_ (.A(_14327_),
    .ZN(_14330_));
 OR4_X1 _31908_ (.A1(\g_row[1].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08265_));
 OAI21_X2 _31909_ (.A(_07394_),
    .B1(_08265_),
    .B2(\g_row[1].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08266_));
 AND4_X1 _31910_ (.A1(\g_row[1].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08267_));
 AOI21_X4 _31911_ (.A(_07398_),
    .B1(_08267_),
    .B2(\g_row[1].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08268_));
 INV_X1 _31912_ (.A(_14329_),
    .ZN(_08269_));
 AOI21_X1 _31913_ (.A(_08266_),
    .B1(_08268_),
    .B2(_08269_),
    .ZN(_00289_));
 INV_X1 _31914_ (.A(_19826_),
    .ZN(_08270_));
 AOI21_X1 _31915_ (.A(_08266_),
    .B1(_08268_),
    .B2(_08270_),
    .ZN(_00290_));
 INV_X1 _31916_ (.A(_14337_),
    .ZN(_08271_));
 AOI21_X1 _31917_ (.A(_08266_),
    .B1(_08268_),
    .B2(_08271_),
    .ZN(_00291_));
 XOR2_X1 _31918_ (.A(_14336_),
    .B(_19835_),
    .Z(_08272_));
 AOI21_X1 _31919_ (.A(_08266_),
    .B1(_08268_),
    .B2(_08272_),
    .ZN(_00292_));
 AOI21_X1 _31920_ (.A(_19830_),
    .B1(_19831_),
    .B2(_19825_),
    .ZN(_08273_));
 INV_X1 _31921_ (.A(_08273_),
    .ZN(_08274_));
 AOI21_X1 _31922_ (.A(_19834_),
    .B1(_08274_),
    .B2(_19835_),
    .ZN(_08275_));
 XNOR2_X1 _31923_ (.A(\g_row[1].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_19832_),
    .ZN(_08276_));
 XNOR2_X1 _31924_ (.A(_07392_),
    .B(_08276_),
    .ZN(_08277_));
 XNOR2_X1 _31925_ (.A(_08275_),
    .B(_08277_),
    .ZN(_08278_));
 AOI21_X1 _31926_ (.A(_08266_),
    .B1(_08268_),
    .B2(_08278_),
    .ZN(_00293_));
 INV_X1 _31927_ (.A(_08266_),
    .ZN(_08279_));
 NAND2_X1 _31928_ (.A1(_08279_),
    .A2(_08268_),
    .ZN(_08280_));
 CLKBUF_X3 _31929_ (.A(_08280_),
    .Z(_08281_));
 NAND2_X1 _31930_ (.A1(_08211_),
    .A2(_08150_),
    .ZN(_08282_));
 INV_X1 _31931_ (.A(_19839_),
    .ZN(_08283_));
 MUX2_X1 _31932_ (.A(_08282_),
    .B(_08283_),
    .S(_14327_),
    .Z(_08284_));
 NOR2_X1 _31933_ (.A1(_08281_),
    .A2(_08284_),
    .ZN(_00288_));
 XOR2_X1 _31934_ (.A(_19838_),
    .B(_08210_),
    .Z(_08285_));
 MUX2_X1 _31935_ (.A(_08283_),
    .B(_08285_),
    .S(_14327_),
    .Z(_08286_));
 NOR2_X1 _31936_ (.A1(_08281_),
    .A2(_08286_),
    .ZN(_00294_));
 NOR2_X1 _31937_ (.A1(_08281_),
    .A2(_08285_),
    .ZN(_08287_));
 XNOR2_X1 _31938_ (.A(_08213_),
    .B(_08217_),
    .ZN(_08288_));
 NOR2_X1 _31939_ (.A1(_08281_),
    .A2(_08288_),
    .ZN(_08289_));
 MUX2_X1 _31940_ (.A(_08287_),
    .B(_08289_),
    .S(_14327_),
    .Z(_00295_));
 NAND2_X1 _31941_ (.A1(_19838_),
    .A2(_08217_),
    .ZN(_08290_));
 NOR2_X1 _31942_ (.A1(_08210_),
    .A2(_08290_),
    .ZN(_08291_));
 XNOR2_X1 _31943_ (.A(_08209_),
    .B(_08291_),
    .ZN(_08292_));
 NOR2_X1 _31944_ (.A1(_08281_),
    .A2(_08292_),
    .ZN(_08293_));
 MUX2_X1 _31945_ (.A(_08289_),
    .B(_08293_),
    .S(_14327_),
    .Z(_00296_));
 XNOR2_X1 _31946_ (.A(_08218_),
    .B(_08223_),
    .ZN(_08294_));
 NOR2_X1 _31947_ (.A1(_08281_),
    .A2(_08294_),
    .ZN(_08295_));
 MUX2_X1 _31948_ (.A(_08293_),
    .B(_08295_),
    .S(_14327_),
    .Z(_00297_));
 INV_X1 _31949_ (.A(_08228_),
    .ZN(_08296_));
 NAND3_X1 _31950_ (.A1(_08209_),
    .A2(_08223_),
    .A3(_08291_),
    .ZN(_08297_));
 XNOR2_X1 _31951_ (.A(_08296_),
    .B(_08297_),
    .ZN(_08298_));
 NOR2_X1 _31952_ (.A1(_08281_),
    .A2(_08298_),
    .ZN(_08299_));
 MUX2_X1 _31953_ (.A(_08295_),
    .B(_08299_),
    .S(_14327_),
    .Z(_00298_));
 XNOR2_X1 _31954_ (.A(_08229_),
    .B(_08232_),
    .ZN(_08300_));
 NOR2_X1 _31955_ (.A1(_08280_),
    .A2(_08300_),
    .ZN(_08301_));
 MUX2_X1 _31956_ (.A(_08299_),
    .B(_08301_),
    .S(_14327_),
    .Z(_00299_));
 OR3_X1 _31957_ (.A1(_08296_),
    .A2(_08232_),
    .A3(_08297_),
    .ZN(_08302_));
 XNOR2_X1 _31958_ (.A(_08202_),
    .B(_08302_),
    .ZN(_08303_));
 NOR2_X1 _31959_ (.A1(_08281_),
    .A2(_08303_),
    .ZN(_08304_));
 MUX2_X1 _31960_ (.A(_08301_),
    .B(_08304_),
    .S(_14327_),
    .Z(_00300_));
 INV_X1 _31961_ (.A(_08262_),
    .ZN(_08305_));
 AND3_X1 _31962_ (.A1(_08233_),
    .A2(_08305_),
    .A3(_08303_),
    .ZN(_08306_));
 AOI21_X1 _31963_ (.A(_08303_),
    .B1(_08263_),
    .B2(_08233_),
    .ZN(_08307_));
 NOR2_X1 _31964_ (.A1(_08179_),
    .A2(_08307_),
    .ZN(_08308_));
 INV_X1 _31965_ (.A(_08178_),
    .ZN(_08309_));
 AOI21_X2 _31966_ (.A(_19783_),
    .B1(_19784_),
    .B2(_08309_),
    .ZN(_08310_));
 OR2_X1 _31967_ (.A1(_08233_),
    .A2(_08305_),
    .ZN(_08311_));
 NAND3_X1 _31968_ (.A1(_08233_),
    .A2(_08250_),
    .A3(_08305_),
    .ZN(_08312_));
 AOI21_X1 _31969_ (.A(_08310_),
    .B1(_08311_),
    .B2(_08312_),
    .ZN(_08313_));
 NOR4_X1 _31970_ (.A1(_08281_),
    .A2(_08306_),
    .A3(_08308_),
    .A4(_08313_),
    .ZN(_00301_));
 NOR2_X1 _31971_ (.A1(_08202_),
    .A2(_08302_),
    .ZN(_08314_));
 OR4_X1 _31972_ (.A1(_08310_),
    .A2(_08233_),
    .A3(_08250_),
    .A4(_08314_),
    .ZN(_08315_));
 AND3_X1 _31973_ (.A1(_08179_),
    .A2(_08250_),
    .A3(_08314_),
    .ZN(_08316_));
 OAI21_X1 _31974_ (.A(_08233_),
    .B1(_08250_),
    .B2(_08314_),
    .ZN(_08317_));
 AOI21_X1 _31975_ (.A(_08316_),
    .B1(_08317_),
    .B2(_08310_),
    .ZN(_08318_));
 NOR2_X1 _31976_ (.A1(_08310_),
    .A2(_08250_),
    .ZN(_08319_));
 AOI21_X1 _31977_ (.A(_08319_),
    .B1(_08233_),
    .B2(_08310_),
    .ZN(_08320_));
 MUX2_X1 _31978_ (.A(_08318_),
    .B(_08320_),
    .S(_08262_),
    .Z(_08321_));
 AOI21_X1 _31979_ (.A(_08281_),
    .B1(_08315_),
    .B2(_08321_),
    .ZN(_00302_));
 CLKBUF_X2 _31980_ (.A(_19863_),
    .Z(_08322_));
 AOI21_X1 _31981_ (.A(_19862_),
    .B1(_08322_),
    .B2(_19864_),
    .ZN(_08323_));
 BUF_X1 _31982_ (.A(_19865_),
    .Z(_08324_));
 NAND2_X1 _31983_ (.A1(_08322_),
    .A2(_08324_),
    .ZN(_08325_));
 CLKBUF_X2 _31984_ (.A(_19868_),
    .Z(_08326_));
 AOI21_X1 _31985_ (.A(_19866_),
    .B1(_19867_),
    .B2(_08326_),
    .ZN(_08327_));
 OAI21_X1 _31986_ (.A(_08323_),
    .B1(_08325_),
    .B2(_08327_),
    .ZN(_08328_));
 INV_X1 _31987_ (.A(_19870_),
    .ZN(_08329_));
 CLKBUF_X2 _31988_ (.A(_19872_),
    .Z(_08330_));
 INV_X1 _31989_ (.A(_19874_),
    .ZN(_08331_));
 AOI21_X1 _31990_ (.A(_19876_),
    .B1(_19877_),
    .B2(_19878_),
    .ZN(_08332_));
 INV_X1 _31991_ (.A(_19875_),
    .ZN(_08333_));
 OAI21_X1 _31992_ (.A(_08331_),
    .B1(_08332_),
    .B2(_08333_),
    .ZN(_08334_));
 CLKBUF_X2 _31993_ (.A(_19873_),
    .Z(_08335_));
 AOI21_X1 _31994_ (.A(_08330_),
    .B1(_08334_),
    .B2(_08335_),
    .ZN(_08336_));
 INV_X1 _31995_ (.A(_19871_),
    .ZN(_08337_));
 OAI21_X2 _31996_ (.A(_08329_),
    .B1(_08336_),
    .B2(_08337_),
    .ZN(_08338_));
 INV_X1 _31997_ (.A(_19867_),
    .ZN(_08339_));
 CLKBUF_X2 _31998_ (.A(_19869_),
    .Z(_08340_));
 INV_X1 _31999_ (.A(_08340_),
    .ZN(_08341_));
 NOR3_X2 _32000_ (.A1(_08339_),
    .A2(_08341_),
    .A3(_08325_),
    .ZN(_08342_));
 AOI21_X2 _32001_ (.A(_08328_),
    .B1(_08338_),
    .B2(_08342_),
    .ZN(_08343_));
 XNOR2_X2 _32002_ (.A(_19861_),
    .B(_08343_),
    .ZN(_08344_));
 INV_X1 _32003_ (.A(_08344_),
    .ZN(_08345_));
 INV_X1 _32004_ (.A(_19866_),
    .ZN(_08346_));
 AOI21_X1 _32005_ (.A(_08326_),
    .B1(_08340_),
    .B2(_08338_),
    .ZN(_08347_));
 OAI21_X2 _32006_ (.A(_08346_),
    .B1(_08347_),
    .B2(_08339_),
    .ZN(_08348_));
 XNOR2_X1 _32007_ (.A(_08324_),
    .B(_08348_),
    .ZN(_08349_));
 XNOR2_X1 _32008_ (.A(_08341_),
    .B(_08338_),
    .ZN(_08350_));
 INV_X1 _32009_ (.A(_19860_),
    .ZN(_08351_));
 INV_X1 _32010_ (.A(_19861_),
    .ZN(_08352_));
 AOI21_X1 _32011_ (.A(_19864_),
    .B1(_08324_),
    .B2(_19866_),
    .ZN(_08353_));
 INV_X1 _32012_ (.A(_08353_),
    .ZN(_08354_));
 AOI21_X1 _32013_ (.A(_19862_),
    .B1(_08354_),
    .B2(_08322_),
    .ZN(_08355_));
 OAI21_X1 _32014_ (.A(_08351_),
    .B1(_08352_),
    .B2(_08355_),
    .ZN(_08356_));
 INV_X1 _32015_ (.A(_08322_),
    .ZN(_08357_));
 NAND2_X1 _32016_ (.A1(_08324_),
    .A2(_19867_),
    .ZN(_08358_));
 NOR3_X2 _32017_ (.A1(_08352_),
    .A2(_08357_),
    .A3(_08358_),
    .ZN(_08359_));
 AOI21_X2 _32018_ (.A(_08326_),
    .B1(_08340_),
    .B2(_19870_),
    .ZN(_08360_));
 OAI21_X1 _32019_ (.A(_08331_),
    .B1(_08333_),
    .B2(_14341_),
    .ZN(_08361_));
 AOI21_X1 _32020_ (.A(_08330_),
    .B1(_08361_),
    .B2(_08335_),
    .ZN(_08362_));
 NAND2_X1 _32021_ (.A1(_08340_),
    .A2(_19871_),
    .ZN(_08363_));
 NOR2_X1 _32022_ (.A1(_08362_),
    .A2(_08363_),
    .ZN(_08364_));
 INV_X1 _32023_ (.A(_08364_),
    .ZN(_08365_));
 NAND2_X1 _32024_ (.A1(_08360_),
    .A2(_08365_),
    .ZN(_08366_));
 AOI21_X1 _32025_ (.A(_08356_),
    .B1(_08359_),
    .B2(_08366_),
    .ZN(_08367_));
 XNOR2_X1 _32026_ (.A(_19859_),
    .B(_08367_),
    .ZN(_19893_));
 AOI21_X1 _32027_ (.A(_08341_),
    .B1(_08337_),
    .B2(_08329_),
    .ZN(_08368_));
 NOR2_X1 _32028_ (.A1(_08326_),
    .A2(_08368_),
    .ZN(_08369_));
 XNOR2_X1 _32029_ (.A(_08339_),
    .B(_08369_),
    .ZN(_08370_));
 XNOR2_X1 _32030_ (.A(_14341_),
    .B(_19875_),
    .ZN(_08371_));
 NOR4_X2 _32031_ (.A1(_14342_),
    .A2(\g_row[1].g_col[3].mult.adder.a[0] ),
    .A3(_19879_),
    .A4(_08371_),
    .ZN(_08372_));
 XNOR2_X1 _32032_ (.A(_08337_),
    .B(_08362_),
    .ZN(_08373_));
 XNOR2_X1 _32033_ (.A(_08335_),
    .B(_08334_),
    .ZN(_08374_));
 NAND4_X1 _32034_ (.A1(_08370_),
    .A2(_08372_),
    .A3(_08373_),
    .A4(_08374_),
    .ZN(_08375_));
 OAI21_X1 _32035_ (.A(_08353_),
    .B1(_08358_),
    .B2(_08360_),
    .ZN(_08376_));
 NOR2_X1 _32036_ (.A1(_08358_),
    .A2(_08365_),
    .ZN(_08377_));
 NOR2_X1 _32037_ (.A1(_08376_),
    .A2(_08377_),
    .ZN(_08378_));
 XNOR2_X1 _32038_ (.A(_08322_),
    .B(_08378_),
    .ZN(_08379_));
 NOR4_X1 _32039_ (.A1(_08350_),
    .A2(_19893_),
    .A3(_08375_),
    .A4(_08379_),
    .ZN(_08380_));
 AND2_X2 _32040_ (.A1(_08349_),
    .A2(_08380_),
    .ZN(_08381_));
 NOR2_X1 _32041_ (.A1(_08345_),
    .A2(_08381_),
    .ZN(_19894_));
 INV_X1 _32042_ (.A(_19840_),
    .ZN(_08382_));
 INV_X1 _32043_ (.A(_19841_),
    .ZN(_08383_));
 BUF_X2 _32044_ (.A(_19843_),
    .Z(_08384_));
 INV_X1 _32045_ (.A(_19844_),
    .ZN(_08385_));
 INV_X1 _32046_ (.A(_19845_),
    .ZN(_08386_));
 INV_X1 _32047_ (.A(_19850_),
    .ZN(_08387_));
 BUF_X2 _32048_ (.A(_19853_),
    .Z(_08388_));
 AOI21_X2 _32049_ (.A(_19852_),
    .B1(_08388_),
    .B2(_19854_),
    .ZN(_08389_));
 CLKBUF_X2 _32050_ (.A(_19851_),
    .Z(_08390_));
 INV_X1 _32051_ (.A(_08390_),
    .ZN(_08391_));
 OAI21_X1 _32052_ (.A(_08387_),
    .B1(_08389_),
    .B2(_08391_),
    .ZN(_08392_));
 AOI21_X1 _32053_ (.A(_19848_),
    .B1(_19849_),
    .B2(_08392_),
    .ZN(_08393_));
 BUF_X2 _32054_ (.A(_19857_),
    .Z(_08394_));
 AND2_X1 _32055_ (.A1(_08394_),
    .A2(_19859_),
    .ZN(_08395_));
 AOI21_X1 _32056_ (.A(_19862_),
    .B1(_08376_),
    .B2(_08322_),
    .ZN(_08396_));
 OAI21_X1 _32057_ (.A(_08351_),
    .B1(_08352_),
    .B2(_08396_),
    .ZN(_08397_));
 AOI221_X2 _32058_ (.A(_19856_),
    .B1(_08394_),
    .B2(_19858_),
    .C1(_08395_),
    .C2(_08397_),
    .ZN(_08398_));
 BUF_X2 _32059_ (.A(_19855_),
    .Z(_08399_));
 NAND4_X1 _32060_ (.A1(_19849_),
    .A2(_08390_),
    .A3(_08388_),
    .A4(_08399_),
    .ZN(_08400_));
 OAI21_X1 _32061_ (.A(_08393_),
    .B1(_08398_),
    .B2(_08400_),
    .ZN(_08401_));
 CLKBUF_X2 _32062_ (.A(_19847_),
    .Z(_08402_));
 AOI21_X1 _32063_ (.A(_19846_),
    .B1(_08401_),
    .B2(_08402_),
    .ZN(_08403_));
 OAI21_X1 _32064_ (.A(_08385_),
    .B1(_08386_),
    .B2(_08403_),
    .ZN(_08404_));
 AOI21_X2 _32065_ (.A(_19842_),
    .B1(_08384_),
    .B2(_08404_),
    .ZN(_08405_));
 OAI21_X4 _32066_ (.A(_08382_),
    .B1(_08383_),
    .B2(_08405_),
    .ZN(_08406_));
 INV_X1 _32067_ (.A(_19852_),
    .ZN(_08407_));
 INV_X1 _32068_ (.A(_08388_),
    .ZN(_08408_));
 AOI21_X1 _32069_ (.A(_19854_),
    .B1(_08399_),
    .B2(_19856_),
    .ZN(_08409_));
 OAI21_X1 _32070_ (.A(_08407_),
    .B1(_08408_),
    .B2(_08409_),
    .ZN(_08410_));
 AOI21_X1 _32071_ (.A(_19850_),
    .B1(_08410_),
    .B2(_08390_),
    .ZN(_08411_));
 NAND4_X1 _32072_ (.A1(_08390_),
    .A2(_08388_),
    .A3(_08399_),
    .A4(_08394_),
    .ZN(_08412_));
 AOI21_X1 _32073_ (.A(_19858_),
    .B1(_19859_),
    .B2(_19860_),
    .ZN(_08413_));
 NAND2_X1 _32074_ (.A1(_19859_),
    .A2(_19861_),
    .ZN(_08414_));
 OAI21_X1 _32075_ (.A(_08413_),
    .B1(_08414_),
    .B2(_08323_),
    .ZN(_08415_));
 NOR2_X1 _32076_ (.A1(_08325_),
    .A2(_08414_),
    .ZN(_08416_));
 INV_X1 _32077_ (.A(_08330_),
    .ZN(_08417_));
 OAI21_X1 _32078_ (.A(_08329_),
    .B1(_08417_),
    .B2(_08337_),
    .ZN(_08418_));
 AOI21_X1 _32079_ (.A(_08326_),
    .B1(_08340_),
    .B2(_08418_),
    .ZN(_08419_));
 OAI21_X1 _32080_ (.A(_08346_),
    .B1(_08419_),
    .B2(_08339_),
    .ZN(_08420_));
 AOI21_X1 _32081_ (.A(_08415_),
    .B1(_08416_),
    .B2(_08420_),
    .ZN(_08421_));
 OAI21_X1 _32082_ (.A(_08411_),
    .B1(_08412_),
    .B2(_08421_),
    .ZN(_08422_));
 AOI21_X1 _32083_ (.A(_19848_),
    .B1(_19849_),
    .B2(_08422_),
    .ZN(_08423_));
 INV_X1 _32084_ (.A(_08423_),
    .ZN(_08424_));
 AOI21_X1 _32085_ (.A(_19846_),
    .B1(_08424_),
    .B2(_08402_),
    .ZN(_08425_));
 OAI21_X1 _32086_ (.A(_08385_),
    .B1(_08386_),
    .B2(_08425_),
    .ZN(_08426_));
 AOI21_X1 _32087_ (.A(_19842_),
    .B1(_08384_),
    .B2(_08426_),
    .ZN(_08427_));
 XNOR2_X1 _32088_ (.A(_19841_),
    .B(_08427_),
    .ZN(_08428_));
 INV_X1 _32089_ (.A(_08428_),
    .ZN(_08429_));
 INV_X1 _32090_ (.A(_19848_),
    .ZN(_08430_));
 INV_X1 _32091_ (.A(_19849_),
    .ZN(_08431_));
 AOI21_X2 _32092_ (.A(_19856_),
    .B1(_08394_),
    .B2(_19858_),
    .ZN(_08432_));
 NAND2_X1 _32093_ (.A1(_08388_),
    .A2(_08399_),
    .ZN(_08433_));
 NAND3_X1 _32094_ (.A1(_08388_),
    .A2(_08399_),
    .A3(_08395_),
    .ZN(_08434_));
 AOI21_X1 _32095_ (.A(_08330_),
    .B1(_19874_),
    .B2(_08335_),
    .ZN(_08435_));
 OAI21_X1 _32096_ (.A(_08360_),
    .B1(_08363_),
    .B2(_08435_),
    .ZN(_08436_));
 AOI21_X1 _32097_ (.A(_08356_),
    .B1(_08359_),
    .B2(_08436_),
    .ZN(_08437_));
 OAI221_X1 _32098_ (.A(_08389_),
    .B1(_08432_),
    .B2(_08433_),
    .C1(_08434_),
    .C2(_08437_),
    .ZN(_08438_));
 AOI21_X1 _32099_ (.A(_19850_),
    .B1(_08438_),
    .B2(_08390_),
    .ZN(_08439_));
 OAI21_X1 _32100_ (.A(_08430_),
    .B1(_08431_),
    .B2(_08439_),
    .ZN(_08440_));
 AOI21_X1 _32101_ (.A(_19846_),
    .B1(_08440_),
    .B2(_08402_),
    .ZN(_08441_));
 OAI21_X2 _32102_ (.A(_08385_),
    .B1(_08386_),
    .B2(_08441_),
    .ZN(_08442_));
 XNOR2_X2 _32103_ (.A(_08384_),
    .B(_08442_),
    .ZN(_08443_));
 NAND2_X1 _32104_ (.A1(_08359_),
    .A2(_08395_),
    .ZN(_08444_));
 OAI21_X2 _32105_ (.A(_08398_),
    .B1(_08444_),
    .B2(_08365_),
    .ZN(_08445_));
 INV_X1 _32106_ (.A(_08445_),
    .ZN(_08446_));
 OAI21_X1 _32107_ (.A(_08393_),
    .B1(_08400_),
    .B2(_08446_),
    .ZN(_08447_));
 XOR2_X2 _32108_ (.A(_08402_),
    .B(_08447_),
    .Z(_08448_));
 NAND2_X1 _32109_ (.A1(_08399_),
    .A2(_08394_),
    .ZN(_08449_));
 OAI21_X1 _32110_ (.A(_08409_),
    .B1(_08449_),
    .B2(_08413_),
    .ZN(_08450_));
 INV_X1 _32111_ (.A(_19876_),
    .ZN(_08451_));
 OAI21_X1 _32112_ (.A(_08331_),
    .B1(_08451_),
    .B2(_08333_),
    .ZN(_08452_));
 AOI21_X1 _32113_ (.A(_08330_),
    .B1(_08452_),
    .B2(_08335_),
    .ZN(_08453_));
 OAI21_X1 _32114_ (.A(_08329_),
    .B1(_08453_),
    .B2(_08337_),
    .ZN(_08454_));
 AOI21_X1 _32115_ (.A(_08328_),
    .B1(_08342_),
    .B2(_08454_),
    .ZN(_08455_));
 NOR3_X1 _32116_ (.A1(_08449_),
    .A2(_08414_),
    .A3(_08455_),
    .ZN(_08456_));
 OAI21_X1 _32117_ (.A(_08388_),
    .B1(_08450_),
    .B2(_08456_),
    .ZN(_08457_));
 NAND2_X1 _32118_ (.A1(_08407_),
    .A2(_08457_),
    .ZN(_08458_));
 AOI21_X1 _32119_ (.A(_19850_),
    .B1(_08458_),
    .B2(_08390_),
    .ZN(_08459_));
 OAI21_X1 _32120_ (.A(_08430_),
    .B1(_08431_),
    .B2(_08459_),
    .ZN(_08460_));
 AOI21_X1 _32121_ (.A(_19846_),
    .B1(_08460_),
    .B2(_08402_),
    .ZN(_08461_));
 XNOR2_X1 _32122_ (.A(_19845_),
    .B(_08461_),
    .ZN(_08462_));
 OAI221_X2 _32123_ (.A(_08389_),
    .B1(_08432_),
    .B2(_08433_),
    .C1(_08434_),
    .C2(_08367_),
    .ZN(_08463_));
 XNOR2_X2 _32124_ (.A(_08391_),
    .B(_08463_),
    .ZN(_08464_));
 AOI21_X2 _32125_ (.A(_08415_),
    .B1(_08416_),
    .B2(_08348_),
    .ZN(_08465_));
 XNOR2_X2 _32126_ (.A(_08394_),
    .B(_08465_),
    .ZN(_08466_));
 AND3_X1 _32127_ (.A1(_08344_),
    .A2(_19893_),
    .A3(_08466_),
    .ZN(_08467_));
 NOR3_X1 _32128_ (.A1(_08343_),
    .A2(_08449_),
    .A3(_08414_),
    .ZN(_08468_));
 NOR2_X1 _32129_ (.A1(_08450_),
    .A2(_08468_),
    .ZN(_08469_));
 XNOR2_X2 _32130_ (.A(_08408_),
    .B(_08469_),
    .ZN(_08470_));
 INV_X1 _32131_ (.A(_08470_),
    .ZN(_08471_));
 XOR2_X2 _32132_ (.A(_08399_),
    .B(_08445_),
    .Z(_08472_));
 AND3_X1 _32133_ (.A1(_08467_),
    .A2(_08471_),
    .A3(_08472_),
    .ZN(_08473_));
 OAI21_X1 _32134_ (.A(_08411_),
    .B1(_08412_),
    .B2(_08465_),
    .ZN(_08474_));
 XNOR2_X2 _32135_ (.A(_08431_),
    .B(_08474_),
    .ZN(_08475_));
 NAND3_X1 _32136_ (.A1(_08464_),
    .A2(_08473_),
    .A3(_08475_),
    .ZN(_08476_));
 INV_X1 _32137_ (.A(_08476_),
    .ZN(_08477_));
 NAND3_X1 _32138_ (.A1(_08448_),
    .A2(_08462_),
    .A3(_08477_),
    .ZN(_08478_));
 NOR3_X1 _32139_ (.A1(_08429_),
    .A2(_08443_),
    .A3(_08478_),
    .ZN(_08479_));
 XOR2_X1 _32140_ (.A(_08406_),
    .B(_08479_),
    .Z(_14344_));
 INV_X1 _32141_ (.A(_14344_),
    .ZN(_14347_));
 OR4_X1 _32142_ (.A1(\g_row[1].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08480_));
 OAI21_X2 _32143_ (.A(_07621_),
    .B1(_08480_),
    .B2(\g_row[1].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08481_));
 AND4_X1 _32144_ (.A1(\g_row[1].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[1].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[1].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[1].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08482_));
 AOI21_X4 _32145_ (.A(_07625_),
    .B1(_08482_),
    .B2(\g_row[1].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08483_));
 INV_X1 _32146_ (.A(_14346_),
    .ZN(_08484_));
 AOI21_X1 _32147_ (.A(_08481_),
    .B1(_08483_),
    .B2(_08484_),
    .ZN(_00305_));
 INV_X1 _32148_ (.A(_19883_),
    .ZN(_08485_));
 AOI21_X1 _32149_ (.A(_08481_),
    .B1(_08483_),
    .B2(_08485_),
    .ZN(_00306_));
 INV_X1 _32150_ (.A(_14354_),
    .ZN(_08486_));
 AOI21_X1 _32151_ (.A(_08481_),
    .B1(_08483_),
    .B2(_08486_),
    .ZN(_00307_));
 XOR2_X1 _32152_ (.A(_14353_),
    .B(_19892_),
    .Z(_08487_));
 AOI21_X1 _32153_ (.A(_08481_),
    .B1(_08483_),
    .B2(_08487_),
    .ZN(_00308_));
 AOI21_X1 _32154_ (.A(_19887_),
    .B1(_19888_),
    .B2(_19882_),
    .ZN(_08488_));
 INV_X1 _32155_ (.A(_08488_),
    .ZN(_08489_));
 AOI21_X1 _32156_ (.A(_19891_),
    .B1(_08489_),
    .B2(_19892_),
    .ZN(_08490_));
 XNOR2_X1 _32157_ (.A(\g_row[1].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_19889_),
    .ZN(_08491_));
 XNOR2_X1 _32158_ (.A(_07619_),
    .B(_08491_),
    .ZN(_08492_));
 XNOR2_X1 _32159_ (.A(_08490_),
    .B(_08492_),
    .ZN(_08493_));
 AOI21_X1 _32160_ (.A(_08481_),
    .B1(_08483_),
    .B2(_08493_),
    .ZN(_00309_));
 INV_X1 _32161_ (.A(_08481_),
    .ZN(_08494_));
 NAND2_X2 _32162_ (.A1(_08494_),
    .A2(_08483_),
    .ZN(_08495_));
 NAND2_X1 _32163_ (.A1(_19896_),
    .A2(_14344_),
    .ZN(_08496_));
 NAND3_X1 _32164_ (.A1(_08344_),
    .A2(_08381_),
    .A3(_14347_),
    .ZN(_08497_));
 AOI21_X1 _32165_ (.A(_08495_),
    .B1(_08496_),
    .B2(_08497_),
    .ZN(_00304_));
 INV_X1 _32166_ (.A(_19896_),
    .ZN(_08498_));
 XNOR2_X2 _32167_ (.A(_19895_),
    .B(_08466_),
    .ZN(_08499_));
 MUX2_X1 _32168_ (.A(_08498_),
    .B(_08499_),
    .S(_14344_),
    .Z(_08500_));
 NOR2_X1 _32169_ (.A1(_08495_),
    .A2(_08500_),
    .ZN(_00310_));
 XNOR2_X1 _32170_ (.A(_08467_),
    .B(_08472_),
    .ZN(_08501_));
 MUX2_X2 _32171_ (.A(_08499_),
    .B(_08501_),
    .S(_14344_),
    .Z(_08502_));
 NOR2_X1 _32172_ (.A1(_08495_),
    .A2(_08502_),
    .ZN(_00311_));
 NAND3_X1 _32173_ (.A1(_19895_),
    .A2(_08466_),
    .A3(_08472_),
    .ZN(_08503_));
 XNOR2_X1 _32174_ (.A(_08470_),
    .B(_08503_),
    .ZN(_08504_));
 MUX2_X2 _32175_ (.A(_08501_),
    .B(_08504_),
    .S(_14344_),
    .Z(_08505_));
 NOR2_X1 _32176_ (.A1(_08495_),
    .A2(_08505_),
    .ZN(_00312_));
 XNOR2_X1 _32177_ (.A(_08464_),
    .B(_08473_),
    .ZN(_08506_));
 MUX2_X2 _32178_ (.A(_08504_),
    .B(_08506_),
    .S(_14344_),
    .Z(_08507_));
 NOR2_X1 _32179_ (.A1(_08495_),
    .A2(_08507_),
    .ZN(_00313_));
 INV_X1 _32180_ (.A(_08464_),
    .ZN(_08508_));
 NOR3_X1 _32181_ (.A1(_08508_),
    .A2(_08470_),
    .A3(_08503_),
    .ZN(_08509_));
 XNOR2_X1 _32182_ (.A(_08475_),
    .B(_08509_),
    .ZN(_08510_));
 MUX2_X2 _32183_ (.A(_08506_),
    .B(_08510_),
    .S(_14344_),
    .Z(_08511_));
 NOR2_X1 _32184_ (.A1(_08495_),
    .A2(_08511_),
    .ZN(_00314_));
 XOR2_X2 _32185_ (.A(_08448_),
    .B(_08476_),
    .Z(_08512_));
 MUX2_X2 _32186_ (.A(_08510_),
    .B(_08512_),
    .S(_14344_),
    .Z(_08513_));
 NOR2_X1 _32187_ (.A1(_08495_),
    .A2(_08513_),
    .ZN(_00315_));
 INV_X1 _32188_ (.A(_08462_),
    .ZN(_08514_));
 NAND3_X1 _32189_ (.A1(_08448_),
    .A2(_08475_),
    .A3(_08509_),
    .ZN(_08515_));
 XNOR2_X1 _32190_ (.A(_08514_),
    .B(_08515_),
    .ZN(_08516_));
 MUX2_X2 _32191_ (.A(_08512_),
    .B(_08516_),
    .S(_14344_),
    .Z(_08517_));
 NOR2_X1 _32192_ (.A1(_08495_),
    .A2(_08517_),
    .ZN(_00316_));
 AND3_X2 _32193_ (.A1(_08448_),
    .A2(_08462_),
    .A3(_08477_),
    .ZN(_08518_));
 XNOR2_X2 _32194_ (.A(_08518_),
    .B(_08443_),
    .ZN(_08519_));
 XOR2_X2 _32195_ (.A(_08384_),
    .B(_08442_),
    .Z(_08520_));
 NOR2_X1 _32196_ (.A1(_08518_),
    .A2(_08520_),
    .ZN(_08521_));
 NAND2_X1 _32197_ (.A1(_08406_),
    .A2(_08428_),
    .ZN(_08522_));
 OAI22_X2 _32198_ (.A1(_08406_),
    .A2(_08479_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08523_));
 INV_X1 _32199_ (.A(_08516_),
    .ZN(_08524_));
 AOI22_X4 _32200_ (.A1(_08406_),
    .A2(_08519_),
    .B1(_08523_),
    .B2(_08524_),
    .ZN(_08525_));
 NOR2_X1 _32201_ (.A1(_08495_),
    .A2(_08525_),
    .ZN(_00317_));
 NOR2_X1 _32202_ (.A1(_08514_),
    .A2(_08515_),
    .ZN(_08526_));
 NAND4_X1 _32203_ (.A1(_08406_),
    .A2(_08429_),
    .A3(_08520_),
    .A4(_08526_),
    .ZN(_08527_));
 OAI21_X1 _32204_ (.A(_08520_),
    .B1(_08526_),
    .B2(_08518_),
    .ZN(_08528_));
 NOR2_X1 _32205_ (.A1(_08406_),
    .A2(_08526_),
    .ZN(_08529_));
 AOI22_X2 _32206_ (.A1(_08406_),
    .A2(_08528_),
    .B1(_08529_),
    .B2(_08518_),
    .ZN(_08530_));
 XNOR2_X1 _32207_ (.A(_08518_),
    .B(_08520_),
    .ZN(_08531_));
 OAI221_X1 _32208_ (.A(_08527_),
    .B1(_08530_),
    .B2(_08429_),
    .C1(_08406_),
    .C2(_08531_),
    .ZN(_08532_));
 AND3_X1 _32209_ (.A1(_08494_),
    .A2(_08483_),
    .A3(_08532_),
    .ZN(_00318_));
 CLKBUF_X2 _32210_ (.A(_19920_),
    .Z(_08533_));
 AOI21_X1 _32211_ (.A(_19919_),
    .B1(_08533_),
    .B2(_19921_),
    .ZN(_08534_));
 BUF_X1 _32212_ (.A(_19922_),
    .Z(_08535_));
 NAND2_X1 _32213_ (.A1(_08533_),
    .A2(_08535_),
    .ZN(_08536_));
 CLKBUF_X2 _32214_ (.A(_19925_),
    .Z(_08537_));
 AOI21_X1 _32215_ (.A(_19923_),
    .B1(_19924_),
    .B2(_08537_),
    .ZN(_08538_));
 OAI21_X1 _32216_ (.A(_08534_),
    .B1(_08536_),
    .B2(_08538_),
    .ZN(_08539_));
 INV_X1 _32217_ (.A(_19927_),
    .ZN(_08540_));
 CLKBUF_X2 _32218_ (.A(_19929_),
    .Z(_08541_));
 INV_X1 _32219_ (.A(_19931_),
    .ZN(_08542_));
 AOI21_X1 _32220_ (.A(_19933_),
    .B1(_19934_),
    .B2(_19935_),
    .ZN(_08543_));
 INV_X1 _32221_ (.A(_19932_),
    .ZN(_08544_));
 OAI21_X1 _32222_ (.A(_08542_),
    .B1(_08543_),
    .B2(_08544_),
    .ZN(_08545_));
 CLKBUF_X2 _32223_ (.A(_19930_),
    .Z(_08546_));
 AOI21_X1 _32224_ (.A(_08541_),
    .B1(_08545_),
    .B2(_08546_),
    .ZN(_08547_));
 INV_X1 _32225_ (.A(_19928_),
    .ZN(_08548_));
 OAI21_X1 _32226_ (.A(_08540_),
    .B1(_08547_),
    .B2(_08548_),
    .ZN(_08549_));
 INV_X1 _32227_ (.A(_19924_),
    .ZN(_08550_));
 CLKBUF_X2 _32228_ (.A(_19926_),
    .Z(_08551_));
 INV_X1 _32229_ (.A(_08551_),
    .ZN(_08552_));
 NOR3_X2 _32230_ (.A1(_08550_),
    .A2(_08552_),
    .A3(_08536_),
    .ZN(_08553_));
 AOI21_X2 _32231_ (.A(_08539_),
    .B1(_08549_),
    .B2(_08553_),
    .ZN(_08554_));
 XNOR2_X1 _32232_ (.A(_19918_),
    .B(_08554_),
    .ZN(_08555_));
 INV_X1 _32233_ (.A(_08555_),
    .ZN(_08556_));
 INV_X1 _32234_ (.A(_19923_),
    .ZN(_08557_));
 AOI21_X1 _32235_ (.A(_08537_),
    .B1(_08551_),
    .B2(_08549_),
    .ZN(_08558_));
 OAI21_X1 _32236_ (.A(_08557_),
    .B1(_08558_),
    .B2(_08550_),
    .ZN(_08559_));
 XNOR2_X1 _32237_ (.A(_08535_),
    .B(_08559_),
    .ZN(_08560_));
 XNOR2_X1 _32238_ (.A(_08552_),
    .B(_08549_),
    .ZN(_08561_));
 INV_X1 _32239_ (.A(_19917_),
    .ZN(_08562_));
 INV_X1 _32240_ (.A(_19918_),
    .ZN(_08563_));
 AOI21_X1 _32241_ (.A(_19921_),
    .B1(_08535_),
    .B2(_19923_),
    .ZN(_08564_));
 INV_X1 _32242_ (.A(_08564_),
    .ZN(_08565_));
 AOI21_X1 _32243_ (.A(_19919_),
    .B1(_08565_),
    .B2(_08533_),
    .ZN(_08566_));
 OAI21_X1 _32244_ (.A(_08562_),
    .B1(_08563_),
    .B2(_08566_),
    .ZN(_08567_));
 INV_X1 _32245_ (.A(_08533_),
    .ZN(_08568_));
 NAND2_X1 _32246_ (.A1(_08535_),
    .A2(_19924_),
    .ZN(_08569_));
 NOR3_X2 _32247_ (.A1(_08563_),
    .A2(_08568_),
    .A3(_08569_),
    .ZN(_08570_));
 AOI21_X2 _32248_ (.A(_08537_),
    .B1(_08551_),
    .B2(_19927_),
    .ZN(_08571_));
 OAI21_X1 _32249_ (.A(_08542_),
    .B1(_08544_),
    .B2(_14358_),
    .ZN(_08572_));
 AOI21_X2 _32250_ (.A(_08541_),
    .B1(_08572_),
    .B2(_08546_),
    .ZN(_08573_));
 NAND2_X1 _32251_ (.A1(_08551_),
    .A2(_19928_),
    .ZN(_08574_));
 NOR2_X1 _32252_ (.A1(_08573_),
    .A2(_08574_),
    .ZN(_08575_));
 INV_X1 _32253_ (.A(_08575_),
    .ZN(_08576_));
 NAND2_X1 _32254_ (.A1(_08571_),
    .A2(_08576_),
    .ZN(_08577_));
 AOI21_X2 _32255_ (.A(_08567_),
    .B1(_08570_),
    .B2(_08577_),
    .ZN(_08578_));
 XNOR2_X1 _32256_ (.A(_19916_),
    .B(_08578_),
    .ZN(_19950_));
 AOI21_X1 _32257_ (.A(_08552_),
    .B1(_08548_),
    .B2(_08540_),
    .ZN(_08579_));
 NOR2_X1 _32258_ (.A1(_08537_),
    .A2(_08579_),
    .ZN(_08580_));
 XNOR2_X1 _32259_ (.A(_08550_),
    .B(_08580_),
    .ZN(_08581_));
 XNOR2_X1 _32260_ (.A(_14358_),
    .B(_19932_),
    .ZN(_08582_));
 NOR4_X1 _32261_ (.A1(_14359_),
    .A2(\g_row[2].g_col[0].mult.adder.a[0] ),
    .A3(_19936_),
    .A4(_08582_),
    .ZN(_08583_));
 XNOR2_X1 _32262_ (.A(_08548_),
    .B(_08573_),
    .ZN(_08584_));
 XNOR2_X1 _32263_ (.A(_08546_),
    .B(_08545_),
    .ZN(_08585_));
 NAND4_X1 _32264_ (.A1(_08581_),
    .A2(_08583_),
    .A3(_08584_),
    .A4(_08585_),
    .ZN(_08586_));
 OAI21_X1 _32265_ (.A(_08564_),
    .B1(_08569_),
    .B2(_08571_),
    .ZN(_08587_));
 NOR2_X1 _32266_ (.A1(_08569_),
    .A2(_08576_),
    .ZN(_08588_));
 NOR2_X1 _32267_ (.A1(_08587_),
    .A2(_08588_),
    .ZN(_08589_));
 XNOR2_X1 _32268_ (.A(_08533_),
    .B(_08589_),
    .ZN(_08590_));
 NOR4_X1 _32269_ (.A1(_08561_),
    .A2(_19950_),
    .A3(_08586_),
    .A4(_08590_),
    .ZN(_08591_));
 AND2_X1 _32270_ (.A1(_08560_),
    .A2(_08591_),
    .ZN(_08592_));
 NOR2_X1 _32271_ (.A1(_08556_),
    .A2(_08592_),
    .ZN(_19951_));
 INV_X1 _32272_ (.A(_19897_),
    .ZN(_08593_));
 INV_X1 _32273_ (.A(_19898_),
    .ZN(_08594_));
 INV_X1 _32274_ (.A(_19901_),
    .ZN(_08595_));
 INV_X1 _32275_ (.A(_19902_),
    .ZN(_08596_));
 CLKBUF_X2 _32276_ (.A(_19906_),
    .Z(_08597_));
 INV_X1 _32277_ (.A(_19907_),
    .ZN(_08598_));
 BUF_X2 _32278_ (.A(_19910_),
    .Z(_08599_));
 AOI21_X2 _32279_ (.A(_19909_),
    .B1(_08599_),
    .B2(_19911_),
    .ZN(_08600_));
 CLKBUF_X2 _32280_ (.A(_19908_),
    .Z(_08601_));
 INV_X1 _32281_ (.A(_08601_),
    .ZN(_08602_));
 OAI21_X1 _32282_ (.A(_08598_),
    .B1(_08600_),
    .B2(_08602_),
    .ZN(_08603_));
 AOI21_X1 _32283_ (.A(_19905_),
    .B1(_08597_),
    .B2(_08603_),
    .ZN(_08604_));
 BUF_X2 _32284_ (.A(_19914_),
    .Z(_08605_));
 AND2_X1 _32285_ (.A1(_08605_),
    .A2(_19916_),
    .ZN(_08606_));
 AOI21_X1 _32286_ (.A(_19919_),
    .B1(_08587_),
    .B2(_08533_),
    .ZN(_08607_));
 OAI21_X1 _32287_ (.A(_08562_),
    .B1(_08563_),
    .B2(_08607_),
    .ZN(_08608_));
 AOI221_X2 _32288_ (.A(_19913_),
    .B1(_08605_),
    .B2(_19915_),
    .C1(_08606_),
    .C2(_08608_),
    .ZN(_08609_));
 BUF_X2 _32289_ (.A(_19912_),
    .Z(_08610_));
 NAND4_X1 _32290_ (.A1(_08597_),
    .A2(_08601_),
    .A3(_08599_),
    .A4(_08610_),
    .ZN(_08611_));
 OAI21_X1 _32291_ (.A(_08604_),
    .B1(_08609_),
    .B2(_08611_),
    .ZN(_08612_));
 CLKBUF_X2 _32292_ (.A(_19904_),
    .Z(_08613_));
 AOI21_X1 _32293_ (.A(_19903_),
    .B1(_08612_),
    .B2(_08613_),
    .ZN(_08614_));
 OAI21_X1 _32294_ (.A(_08595_),
    .B1(_08596_),
    .B2(_08614_),
    .ZN(_08615_));
 AOI21_X1 _32295_ (.A(_19899_),
    .B1(_19900_),
    .B2(_08615_),
    .ZN(_08616_));
 OAI21_X2 _32296_ (.A(_08593_),
    .B1(_08594_),
    .B2(_08616_),
    .ZN(_08617_));
 INV_X1 _32297_ (.A(_19909_),
    .ZN(_08618_));
 INV_X1 _32298_ (.A(_08599_),
    .ZN(_08619_));
 AOI21_X1 _32299_ (.A(_19911_),
    .B1(_08610_),
    .B2(_19913_),
    .ZN(_08620_));
 OAI21_X1 _32300_ (.A(_08618_),
    .B1(_08619_),
    .B2(_08620_),
    .ZN(_08621_));
 AOI21_X1 _32301_ (.A(_19907_),
    .B1(_08621_),
    .B2(_08601_),
    .ZN(_08622_));
 NAND4_X1 _32302_ (.A1(_08601_),
    .A2(_08599_),
    .A3(_08610_),
    .A4(_08605_),
    .ZN(_08623_));
 AOI21_X1 _32303_ (.A(_19915_),
    .B1(_19916_),
    .B2(_19917_),
    .ZN(_08624_));
 NAND2_X1 _32304_ (.A1(_19916_),
    .A2(_19918_),
    .ZN(_08625_));
 OAI21_X1 _32305_ (.A(_08624_),
    .B1(_08625_),
    .B2(_08534_),
    .ZN(_08626_));
 NOR2_X1 _32306_ (.A1(_08536_),
    .A2(_08625_),
    .ZN(_08627_));
 INV_X1 _32307_ (.A(_08541_),
    .ZN(_08628_));
 OAI21_X1 _32308_ (.A(_08540_),
    .B1(_08628_),
    .B2(_08548_),
    .ZN(_08629_));
 AOI21_X1 _32309_ (.A(_08537_),
    .B1(_08551_),
    .B2(_08629_),
    .ZN(_08630_));
 OAI21_X1 _32310_ (.A(_08557_),
    .B1(_08630_),
    .B2(_08550_),
    .ZN(_08631_));
 AOI21_X1 _32311_ (.A(_08626_),
    .B1(_08627_),
    .B2(_08631_),
    .ZN(_08632_));
 OAI21_X1 _32312_ (.A(_08622_),
    .B1(_08623_),
    .B2(_08632_),
    .ZN(_08633_));
 AOI21_X1 _32313_ (.A(_19905_),
    .B1(_08597_),
    .B2(_08633_),
    .ZN(_08634_));
 INV_X1 _32314_ (.A(_08634_),
    .ZN(_08635_));
 AOI21_X1 _32315_ (.A(_19903_),
    .B1(_08635_),
    .B2(_08613_),
    .ZN(_08636_));
 OAI21_X1 _32316_ (.A(_08595_),
    .B1(_08596_),
    .B2(_08636_),
    .ZN(_08637_));
 AOI21_X1 _32317_ (.A(_19899_),
    .B1(_19900_),
    .B2(_08637_),
    .ZN(_08638_));
 XNOR2_X1 _32318_ (.A(_19898_),
    .B(_08638_),
    .ZN(_08639_));
 INV_X1 _32319_ (.A(_08639_),
    .ZN(_08640_));
 INV_X1 _32320_ (.A(_19905_),
    .ZN(_08641_));
 INV_X1 _32321_ (.A(_08597_),
    .ZN(_08642_));
 AOI21_X2 _32322_ (.A(_19913_),
    .B1(_08605_),
    .B2(_19915_),
    .ZN(_08643_));
 NAND2_X1 _32323_ (.A1(_08599_),
    .A2(_08610_),
    .ZN(_08644_));
 NAND3_X1 _32324_ (.A1(_08599_),
    .A2(_08610_),
    .A3(_08606_),
    .ZN(_08645_));
 AOI21_X1 _32325_ (.A(_08541_),
    .B1(_19931_),
    .B2(_08546_),
    .ZN(_08646_));
 OAI21_X1 _32326_ (.A(_08571_),
    .B1(_08574_),
    .B2(_08646_),
    .ZN(_08647_));
 AOI21_X1 _32327_ (.A(_08567_),
    .B1(_08570_),
    .B2(_08647_),
    .ZN(_08648_));
 OAI221_X1 _32328_ (.A(_08600_),
    .B1(_08643_),
    .B2(_08644_),
    .C1(_08645_),
    .C2(_08648_),
    .ZN(_08649_));
 AOI21_X1 _32329_ (.A(_19907_),
    .B1(_08649_),
    .B2(_08601_),
    .ZN(_08650_));
 OAI21_X1 _32330_ (.A(_08641_),
    .B1(_08642_),
    .B2(_08650_),
    .ZN(_08651_));
 AOI21_X1 _32331_ (.A(_19903_),
    .B1(_08651_),
    .B2(_08613_),
    .ZN(_08652_));
 OAI21_X1 _32332_ (.A(_08595_),
    .B1(_08596_),
    .B2(_08652_),
    .ZN(_08653_));
 XOR2_X2 _32333_ (.A(_19900_),
    .B(_08653_),
    .Z(_08654_));
 NAND2_X1 _32334_ (.A1(_08570_),
    .A2(_08606_),
    .ZN(_08655_));
 OAI21_X2 _32335_ (.A(_08609_),
    .B1(_08655_),
    .B2(_08576_),
    .ZN(_08656_));
 INV_X1 _32336_ (.A(_08656_),
    .ZN(_08657_));
 OAI21_X1 _32337_ (.A(_08604_),
    .B1(_08611_),
    .B2(_08657_),
    .ZN(_08658_));
 XNOR2_X2 _32338_ (.A(_08613_),
    .B(_08658_),
    .ZN(_08659_));
 NAND2_X1 _32339_ (.A1(_08610_),
    .A2(_08605_),
    .ZN(_08660_));
 OAI21_X1 _32340_ (.A(_08620_),
    .B1(_08660_),
    .B2(_08624_),
    .ZN(_08661_));
 INV_X1 _32341_ (.A(_19933_),
    .ZN(_08662_));
 OAI21_X1 _32342_ (.A(_08542_),
    .B1(_08662_),
    .B2(_08544_),
    .ZN(_08663_));
 AOI21_X1 _32343_ (.A(_08541_),
    .B1(_08663_),
    .B2(_08546_),
    .ZN(_08664_));
 OAI21_X1 _32344_ (.A(_08540_),
    .B1(_08664_),
    .B2(_08548_),
    .ZN(_08665_));
 AOI21_X1 _32345_ (.A(_08539_),
    .B1(_08553_),
    .B2(_08665_),
    .ZN(_08666_));
 NOR3_X1 _32346_ (.A1(_08660_),
    .A2(_08625_),
    .A3(_08666_),
    .ZN(_08667_));
 OAI21_X1 _32347_ (.A(_08599_),
    .B1(_08661_),
    .B2(_08667_),
    .ZN(_08668_));
 NAND2_X1 _32348_ (.A1(_08618_),
    .A2(_08668_),
    .ZN(_08669_));
 AOI21_X1 _32349_ (.A(_19907_),
    .B1(_08669_),
    .B2(_08601_),
    .ZN(_08670_));
 OAI21_X1 _32350_ (.A(_08641_),
    .B1(_08642_),
    .B2(_08670_),
    .ZN(_08671_));
 AOI21_X1 _32351_ (.A(_19903_),
    .B1(_08671_),
    .B2(_08613_),
    .ZN(_08672_));
 XNOR2_X1 _32352_ (.A(_19902_),
    .B(_08672_),
    .ZN(_08673_));
 INV_X1 _32353_ (.A(_08673_),
    .ZN(_08674_));
 OAI221_X2 _32354_ (.A(_08600_),
    .B1(_08643_),
    .B2(_08644_),
    .C1(_08645_),
    .C2(_08578_),
    .ZN(_08675_));
 XNOR2_X2 _32355_ (.A(_08602_),
    .B(_08675_),
    .ZN(_08676_));
 AOI21_X1 _32356_ (.A(_08626_),
    .B1(_08627_),
    .B2(_08559_),
    .ZN(_08677_));
 XNOR2_X1 _32357_ (.A(_08605_),
    .B(_08677_),
    .ZN(_08678_));
 AND3_X1 _32358_ (.A1(_08555_),
    .A2(_19950_),
    .A3(_08678_),
    .ZN(_08679_));
 NOR3_X1 _32359_ (.A1(_08554_),
    .A2(_08660_),
    .A3(_08625_),
    .ZN(_08680_));
 NOR2_X1 _32360_ (.A1(_08661_),
    .A2(_08680_),
    .ZN(_08681_));
 XNOR2_X1 _32361_ (.A(_08599_),
    .B(_08681_),
    .ZN(_08682_));
 XOR2_X2 _32362_ (.A(_08610_),
    .B(_08656_),
    .Z(_08683_));
 AND3_X1 _32363_ (.A1(_08679_),
    .A2(_08682_),
    .A3(_08683_),
    .ZN(_08684_));
 OAI21_X1 _32364_ (.A(_08622_),
    .B1(_08623_),
    .B2(_08677_),
    .ZN(_08685_));
 XNOR2_X2 _32365_ (.A(_08597_),
    .B(_08685_),
    .ZN(_08686_));
 INV_X1 _32366_ (.A(_08686_),
    .ZN(_08687_));
 NAND3_X1 _32367_ (.A1(_08676_),
    .A2(_08684_),
    .A3(_08687_),
    .ZN(_08688_));
 NOR3_X1 _32368_ (.A1(_08659_),
    .A2(_08674_),
    .A3(_08688_),
    .ZN(_08689_));
 NAND2_X1 _32369_ (.A1(_08654_),
    .A2(_08689_),
    .ZN(_08690_));
 NOR2_X1 _32370_ (.A1(_08640_),
    .A2(_08690_),
    .ZN(_08691_));
 XOR2_X2 _32371_ (.A(_08617_),
    .B(_08691_),
    .Z(_08692_));
 BUF_X1 _32372_ (.A(_08692_),
    .Z(_14361_));
 INV_X1 _32373_ (.A(_14361_),
    .ZN(_14365_));
 OR4_X1 _32374_ (.A1(\g_row[2].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08693_));
 OAI21_X2 _32375_ (.A(_06947_),
    .B1(_08693_),
    .B2(\g_row[2].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08694_));
 AND4_X1 _32376_ (.A1(\g_row[2].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08695_));
 AOI21_X4 _32377_ (.A(_06951_),
    .B1(_08695_),
    .B2(\g_row[2].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08696_));
 INV_X1 _32378_ (.A(_14363_),
    .ZN(_08697_));
 AOI21_X1 _32379_ (.A(_08694_),
    .B1(_08696_),
    .B2(_08697_),
    .ZN(_00321_));
 INV_X1 _32380_ (.A(_19940_),
    .ZN(_08698_));
 AOI21_X1 _32381_ (.A(_08694_),
    .B1(_08696_),
    .B2(_08698_),
    .ZN(_00322_));
 INV_X1 _32382_ (.A(_14371_),
    .ZN(_08699_));
 AOI21_X1 _32383_ (.A(_08694_),
    .B1(_08696_),
    .B2(_08699_),
    .ZN(_00323_));
 XOR2_X1 _32384_ (.A(_14370_),
    .B(_19949_),
    .Z(_08700_));
 AOI21_X1 _32385_ (.A(_08694_),
    .B1(_08696_),
    .B2(_08700_),
    .ZN(_00324_));
 AOI21_X1 _32386_ (.A(_19944_),
    .B1(_19945_),
    .B2(_19939_),
    .ZN(_08701_));
 INV_X1 _32387_ (.A(_08701_),
    .ZN(_08702_));
 AOI21_X1 _32388_ (.A(_19948_),
    .B1(_08702_),
    .B2(_19949_),
    .ZN(_08703_));
 XNOR2_X1 _32389_ (.A(\g_row[2].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_19946_),
    .ZN(_08704_));
 XNOR2_X1 _32390_ (.A(_06945_),
    .B(_08704_),
    .ZN(_08705_));
 XNOR2_X1 _32391_ (.A(_08703_),
    .B(_08705_),
    .ZN(_08706_));
 AOI21_X1 _32392_ (.A(_08694_),
    .B1(_08696_),
    .B2(_08706_),
    .ZN(_00325_));
 INV_X1 _32393_ (.A(_08694_),
    .ZN(_08707_));
 NAND2_X4 _32394_ (.A1(_08707_),
    .A2(_08696_),
    .ZN(_08708_));
 NAND2_X1 _32395_ (.A1(_19953_),
    .A2(_14361_),
    .ZN(_08709_));
 NAND3_X1 _32396_ (.A1(_08555_),
    .A2(_08592_),
    .A3(_14365_),
    .ZN(_08710_));
 AOI21_X1 _32397_ (.A(_08708_),
    .B1(_08709_),
    .B2(_08710_),
    .ZN(_00320_));
 INV_X1 _32398_ (.A(_19953_),
    .ZN(_08711_));
 XNOR2_X1 _32399_ (.A(_19952_),
    .B(_08678_),
    .ZN(_08712_));
 MUX2_X1 _32400_ (.A(_08711_),
    .B(_08712_),
    .S(_14361_),
    .Z(_08713_));
 NOR2_X1 _32401_ (.A1(_08708_),
    .A2(_08713_),
    .ZN(_00326_));
 XNOR2_X1 _32402_ (.A(_08679_),
    .B(_08683_),
    .ZN(_08714_));
 MUX2_X1 _32403_ (.A(_08712_),
    .B(_08714_),
    .S(_14361_),
    .Z(_08715_));
 NOR2_X1 _32404_ (.A1(_08708_),
    .A2(_08715_),
    .ZN(_00327_));
 AND3_X1 _32405_ (.A1(_19952_),
    .A2(_08678_),
    .A3(_08683_),
    .ZN(_08716_));
 XNOR2_X1 _32406_ (.A(_08682_),
    .B(_08716_),
    .ZN(_08717_));
 MUX2_X1 _32407_ (.A(_08714_),
    .B(_08717_),
    .S(_14361_),
    .Z(_08718_));
 NOR2_X1 _32408_ (.A1(_08708_),
    .A2(_08718_),
    .ZN(_00328_));
 XNOR2_X1 _32409_ (.A(_08676_),
    .B(_08684_),
    .ZN(_08719_));
 MUX2_X1 _32410_ (.A(_08717_),
    .B(_08719_),
    .S(_14361_),
    .Z(_08720_));
 NOR2_X1 _32411_ (.A1(_08708_),
    .A2(_08720_),
    .ZN(_00329_));
 AND3_X1 _32412_ (.A1(_08676_),
    .A2(_08682_),
    .A3(_08716_),
    .ZN(_08721_));
 XNOR2_X1 _32413_ (.A(_08687_),
    .B(_08721_),
    .ZN(_08722_));
 MUX2_X1 _32414_ (.A(_08719_),
    .B(_08722_),
    .S(_14361_),
    .Z(_08723_));
 NOR2_X1 _32415_ (.A1(_08708_),
    .A2(_08723_),
    .ZN(_00330_));
 XNOR2_X1 _32416_ (.A(_08659_),
    .B(_08688_),
    .ZN(_08724_));
 MUX2_X1 _32417_ (.A(_08722_),
    .B(_08724_),
    .S(_08692_),
    .Z(_08725_));
 NOR2_X1 _32418_ (.A1(_08708_),
    .A2(_08725_),
    .ZN(_00331_));
 INV_X1 _32419_ (.A(_08721_),
    .ZN(_08726_));
 NOR3_X1 _32420_ (.A1(_08659_),
    .A2(_08686_),
    .A3(_08726_),
    .ZN(_08727_));
 XNOR2_X2 _32421_ (.A(_08674_),
    .B(_08727_),
    .ZN(_08728_));
 NAND2_X1 _32422_ (.A1(_14361_),
    .A2(_08728_),
    .ZN(_08729_));
 OR2_X1 _32423_ (.A1(_14361_),
    .A2(_08724_),
    .ZN(_08730_));
 AOI21_X1 _32424_ (.A(_08708_),
    .B1(_08729_),
    .B2(_08730_),
    .ZN(_00332_));
 NOR2_X1 _32425_ (.A1(_08690_),
    .A2(_08728_),
    .ZN(_08731_));
 OAI21_X1 _32426_ (.A(_08728_),
    .B1(_08690_),
    .B2(_08640_),
    .ZN(_08732_));
 NOR3_X2 _32427_ (.A1(_08659_),
    .A2(_08674_),
    .A3(_08688_),
    .ZN(_08733_));
 OR2_X1 _32428_ (.A1(_08733_),
    .A2(_08654_),
    .ZN(_08734_));
 OAI21_X1 _32429_ (.A(_08734_),
    .B1(_08690_),
    .B2(_08639_),
    .ZN(_08735_));
 MUX2_X1 _32430_ (.A(_08732_),
    .B(_08735_),
    .S(_08617_),
    .Z(_08736_));
 NOR3_X1 _32431_ (.A1(_08708_),
    .A2(_08731_),
    .A3(_08736_),
    .ZN(_00333_));
 AND2_X1 _32432_ (.A1(_08673_),
    .A2(_08727_),
    .ZN(_08737_));
 OAI211_X2 _32433_ (.A(_08733_),
    .B(_08654_),
    .C1(_08737_),
    .C2(_08640_),
    .ZN(_08738_));
 AOI21_X1 _32434_ (.A(_08617_),
    .B1(_08734_),
    .B2(_08738_),
    .ZN(_08739_));
 NAND2_X1 _32435_ (.A1(_08654_),
    .A2(_08737_),
    .ZN(_08740_));
 NAND2_X1 _32436_ (.A1(_08640_),
    .A2(_08740_),
    .ZN(_08741_));
 OAI21_X1 _32437_ (.A(_08654_),
    .B1(_08737_),
    .B2(_08733_),
    .ZN(_08742_));
 OAI21_X1 _32438_ (.A(_08741_),
    .B1(_08742_),
    .B2(_08640_),
    .ZN(_08743_));
 AND2_X1 _32439_ (.A1(_08617_),
    .A2(_08743_),
    .ZN(_08744_));
 NOR3_X1 _32440_ (.A1(_08708_),
    .A2(_08739_),
    .A3(_08744_),
    .ZN(_00334_));
 BUF_X1 _32441_ (.A(_19975_),
    .Z(_08745_));
 INV_X1 _32442_ (.A(_08745_),
    .ZN(_08746_));
 BUF_X1 _32443_ (.A(_19977_),
    .Z(_08747_));
 AOI21_X1 _32444_ (.A(_19976_),
    .B1(_08747_),
    .B2(_19978_),
    .ZN(_08748_));
 BUF_X2 _32445_ (.A(_19979_),
    .Z(_08749_));
 NAND2_X2 _32446_ (.A1(_08747_),
    .A2(_08749_),
    .ZN(_08750_));
 CLKBUF_X2 _32447_ (.A(_19982_),
    .Z(_08751_));
 AOI21_X1 _32448_ (.A(_19980_),
    .B1(_19981_),
    .B2(_08751_),
    .ZN(_08752_));
 OAI21_X1 _32449_ (.A(_08748_),
    .B1(_08750_),
    .B2(_08752_),
    .ZN(_08753_));
 INV_X1 _32450_ (.A(_19984_),
    .ZN(_08754_));
 CLKBUF_X2 _32451_ (.A(_19986_),
    .Z(_08755_));
 INV_X1 _32452_ (.A(_19988_),
    .ZN(_08756_));
 AOI21_X1 _32453_ (.A(_19990_),
    .B1(_19991_),
    .B2(_19992_),
    .ZN(_08757_));
 INV_X1 _32454_ (.A(_19989_),
    .ZN(_08758_));
 OAI21_X1 _32455_ (.A(_08756_),
    .B1(_08757_),
    .B2(_08758_),
    .ZN(_08759_));
 CLKBUF_X2 _32456_ (.A(_19987_),
    .Z(_08760_));
 AOI21_X1 _32457_ (.A(_08755_),
    .B1(_08759_),
    .B2(_08760_),
    .ZN(_08761_));
 INV_X1 _32458_ (.A(_19985_),
    .ZN(_08762_));
 OAI21_X1 _32459_ (.A(_08754_),
    .B1(_08761_),
    .B2(_08762_),
    .ZN(_08763_));
 INV_X2 _32460_ (.A(_19981_),
    .ZN(_08764_));
 CLKBUF_X2 _32461_ (.A(_19983_),
    .Z(_08765_));
 INV_X1 _32462_ (.A(_08765_),
    .ZN(_08766_));
 NOR3_X2 _32463_ (.A1(_08764_),
    .A2(_08766_),
    .A3(_08750_),
    .ZN(_08767_));
 AOI21_X2 _32464_ (.A(_08753_),
    .B1(_08763_),
    .B2(_08767_),
    .ZN(_08768_));
 XNOR2_X1 _32465_ (.A(_08746_),
    .B(_08768_),
    .ZN(_08769_));
 INV_X1 _32466_ (.A(_19980_),
    .ZN(_08770_));
 AOI21_X1 _32467_ (.A(_08751_),
    .B1(_08765_),
    .B2(_08763_),
    .ZN(_08771_));
 OAI21_X1 _32468_ (.A(_08770_),
    .B1(_08771_),
    .B2(_08764_),
    .ZN(_08772_));
 XOR2_X2 _32469_ (.A(_08749_),
    .B(_08772_),
    .Z(_08773_));
 NAND2_X1 _32470_ (.A1(_08764_),
    .A2(_08770_),
    .ZN(_08774_));
 AOI21_X1 _32471_ (.A(_19978_),
    .B1(_08749_),
    .B2(_08774_),
    .ZN(_08775_));
 XNOR2_X1 _32472_ (.A(_08747_),
    .B(_08775_),
    .ZN(_08776_));
 XNOR2_X1 _32473_ (.A(_14375_),
    .B(_19989_),
    .ZN(_08777_));
 OR4_X1 _32474_ (.A1(_14376_),
    .A2(\g_row[2].g_col[1].mult.adder.a[0] ),
    .A3(_19993_),
    .A4(_08777_),
    .ZN(_08778_));
 OAI21_X1 _32475_ (.A(_08756_),
    .B1(_08758_),
    .B2(_14375_),
    .ZN(_08779_));
 AOI21_X2 _32476_ (.A(_08755_),
    .B1(_08779_),
    .B2(_08760_),
    .ZN(_08780_));
 XNOR2_X1 _32477_ (.A(_19985_),
    .B(_08780_),
    .ZN(_08781_));
 NOR3_X1 _32478_ (.A1(_08776_),
    .A2(_08778_),
    .A3(_08781_),
    .ZN(_08782_));
 AOI21_X1 _32479_ (.A(_08766_),
    .B1(_08762_),
    .B2(_08754_),
    .ZN(_08783_));
 NOR2_X1 _32480_ (.A1(_08751_),
    .A2(_08783_),
    .ZN(_08784_));
 XNOR2_X1 _32481_ (.A(_08764_),
    .B(_08784_),
    .ZN(_08785_));
 XNOR2_X1 _32482_ (.A(_08760_),
    .B(_08759_),
    .ZN(_08786_));
 NAND3_X1 _32483_ (.A1(_08782_),
    .A2(_08785_),
    .A3(_08786_),
    .ZN(_08787_));
 CLKBUF_X2 _32484_ (.A(_19973_),
    .Z(_08788_));
 INV_X1 _32485_ (.A(_19976_),
    .ZN(_08789_));
 AOI21_X1 _32486_ (.A(_19978_),
    .B1(_08749_),
    .B2(_19980_),
    .ZN(_08790_));
 INV_X1 _32487_ (.A(_08747_),
    .ZN(_08791_));
 OAI21_X1 _32488_ (.A(_08789_),
    .B1(_08790_),
    .B2(_08791_),
    .ZN(_08792_));
 AND2_X1 _32489_ (.A1(_08745_),
    .A2(_08792_),
    .ZN(_08793_));
 OR2_X1 _32490_ (.A1(_19974_),
    .A2(_08793_),
    .ZN(_08794_));
 NOR3_X2 _32491_ (.A1(_08746_),
    .A2(_08764_),
    .A3(_08750_),
    .ZN(_08795_));
 AOI21_X2 _32492_ (.A(_08751_),
    .B1(_08765_),
    .B2(_19984_),
    .ZN(_08796_));
 NAND2_X1 _32493_ (.A1(_08765_),
    .A2(_19985_),
    .ZN(_08797_));
 OAI21_X1 _32494_ (.A(_08796_),
    .B1(_08797_),
    .B2(_08780_),
    .ZN(_08798_));
 AOI21_X2 _32495_ (.A(_08794_),
    .B1(_08795_),
    .B2(_08798_),
    .ZN(_08799_));
 XNOR2_X2 _32496_ (.A(_08788_),
    .B(_08799_),
    .ZN(_20007_));
 XNOR2_X1 _32497_ (.A(_08766_),
    .B(_08763_),
    .ZN(_08800_));
 NOR4_X1 _32498_ (.A1(_08773_),
    .A2(_08787_),
    .A3(_20007_),
    .A4(_08800_),
    .ZN(_08801_));
 NOR2_X1 _32499_ (.A1(_08769_),
    .A2(_08801_),
    .ZN(_20008_));
 INV_X1 _32500_ (.A(_19956_),
    .ZN(_08802_));
 INV_X1 _32501_ (.A(_19957_),
    .ZN(_08803_));
 BUF_X1 _32502_ (.A(_19959_),
    .Z(_08804_));
 INV_X1 _32503_ (.A(_19960_),
    .ZN(_08805_));
 INV_X1 _32504_ (.A(_19962_),
    .ZN(_08806_));
 INV_X1 _32505_ (.A(_19963_),
    .ZN(_08807_));
 CLKBUF_X2 _32506_ (.A(_19967_),
    .Z(_08808_));
 AOI21_X2 _32507_ (.A(_19966_),
    .B1(_08808_),
    .B2(_19968_),
    .ZN(_08809_));
 INV_X1 _32508_ (.A(_08809_),
    .ZN(_08810_));
 CLKBUF_X2 _32509_ (.A(_19965_),
    .Z(_08811_));
 AOI21_X1 _32510_ (.A(_19964_),
    .B1(_08810_),
    .B2(_08811_),
    .ZN(_08812_));
 OAI21_X1 _32511_ (.A(_08806_),
    .B1(_08807_),
    .B2(_08812_),
    .ZN(_08813_));
 BUF_X2 _32512_ (.A(_19971_),
    .Z(_08814_));
 AOI21_X2 _32513_ (.A(_19970_),
    .B1(_08814_),
    .B2(_19972_),
    .ZN(_08815_));
 NAND2_X1 _32514_ (.A1(_08814_),
    .A2(_08788_),
    .ZN(_08816_));
 OAI21_X1 _32515_ (.A(_08770_),
    .B1(_08796_),
    .B2(_08764_),
    .ZN(_08817_));
 AOI21_X1 _32516_ (.A(_19978_),
    .B1(_08749_),
    .B2(_08817_),
    .ZN(_08818_));
 OAI21_X1 _32517_ (.A(_08789_),
    .B1(_08818_),
    .B2(_08791_),
    .ZN(_08819_));
 AOI21_X1 _32518_ (.A(_19974_),
    .B1(_08745_),
    .B2(_08819_),
    .ZN(_08820_));
 OAI21_X1 _32519_ (.A(_08815_),
    .B1(_08816_),
    .B2(_08820_),
    .ZN(_08821_));
 INV_X1 _32520_ (.A(_08811_),
    .ZN(_08822_));
 BUF_X2 _32521_ (.A(_19969_),
    .Z(_08823_));
 NAND2_X1 _32522_ (.A1(_08808_),
    .A2(_08823_),
    .ZN(_08824_));
 NOR3_X2 _32523_ (.A1(_08807_),
    .A2(_08822_),
    .A3(_08824_),
    .ZN(_08825_));
 AOI21_X1 _32524_ (.A(_08813_),
    .B1(_08821_),
    .B2(_08825_),
    .ZN(_08826_));
 CLKBUF_X2 _32525_ (.A(_19961_),
    .Z(_08827_));
 INV_X1 _32526_ (.A(_08827_),
    .ZN(_08828_));
 OAI21_X1 _32527_ (.A(_08805_),
    .B1(_08826_),
    .B2(_08828_),
    .ZN(_08829_));
 AOI21_X1 _32528_ (.A(_19958_),
    .B1(_08804_),
    .B2(_08829_),
    .ZN(_08830_));
 OAI21_X2 _32529_ (.A(_08802_),
    .B1(_08803_),
    .B2(_08830_),
    .ZN(_08831_));
 AOI21_X4 _32530_ (.A(_19954_),
    .B1(_19955_),
    .B2(_08831_),
    .ZN(_08832_));
 INV_X1 _32531_ (.A(_19966_),
    .ZN(_08833_));
 INV_X1 _32532_ (.A(_08808_),
    .ZN(_08834_));
 AOI21_X1 _32533_ (.A(_19968_),
    .B1(_08823_),
    .B2(_19970_),
    .ZN(_08835_));
 OAI21_X1 _32534_ (.A(_08833_),
    .B1(_08834_),
    .B2(_08835_),
    .ZN(_08836_));
 AOI21_X1 _32535_ (.A(_19964_),
    .B1(_08836_),
    .B2(_08811_),
    .ZN(_08837_));
 NAND4_X1 _32536_ (.A1(_08811_),
    .A2(_08808_),
    .A3(_08823_),
    .A4(_08814_),
    .ZN(_08838_));
 AOI21_X1 _32537_ (.A(_19972_),
    .B1(_08788_),
    .B2(_19974_),
    .ZN(_08839_));
 NAND2_X1 _32538_ (.A1(_08788_),
    .A2(_08745_),
    .ZN(_08840_));
 OAI21_X1 _32539_ (.A(_08839_),
    .B1(_08840_),
    .B2(_08748_),
    .ZN(_08841_));
 NOR2_X1 _32540_ (.A1(_08750_),
    .A2(_08840_),
    .ZN(_08842_));
 INV_X1 _32541_ (.A(_08755_),
    .ZN(_08843_));
 OAI21_X1 _32542_ (.A(_08754_),
    .B1(_08843_),
    .B2(_08762_),
    .ZN(_08844_));
 AOI21_X1 _32543_ (.A(_08751_),
    .B1(_08765_),
    .B2(_08844_),
    .ZN(_08845_));
 OAI21_X1 _32544_ (.A(_08770_),
    .B1(_08845_),
    .B2(_08764_),
    .ZN(_08846_));
 AOI21_X1 _32545_ (.A(_08841_),
    .B1(_08842_),
    .B2(_08846_),
    .ZN(_08847_));
 OAI21_X1 _32546_ (.A(_08837_),
    .B1(_08838_),
    .B2(_08847_),
    .ZN(_08848_));
 AOI21_X1 _32547_ (.A(_19962_),
    .B1(_19963_),
    .B2(_08848_),
    .ZN(_08849_));
 OAI21_X1 _32548_ (.A(_08805_),
    .B1(_08849_),
    .B2(_08828_),
    .ZN(_08850_));
 AOI21_X1 _32549_ (.A(_19958_),
    .B1(_08804_),
    .B2(_08850_),
    .ZN(_08851_));
 OAI21_X1 _32550_ (.A(_08802_),
    .B1(_08803_),
    .B2(_08851_),
    .ZN(_08852_));
 XNOR2_X2 _32551_ (.A(_19955_),
    .B(_08852_),
    .ZN(_08853_));
 NOR4_X1 _32552_ (.A1(_08746_),
    .A2(_08764_),
    .A3(_08750_),
    .A4(_08816_),
    .ZN(_08854_));
 NOR2_X1 _32553_ (.A1(_08780_),
    .A2(_08797_),
    .ZN(_08855_));
 AOI21_X2 _32554_ (.A(_08821_),
    .B1(_08854_),
    .B2(_08855_),
    .ZN(_08856_));
 INV_X1 _32555_ (.A(_08856_),
    .ZN(_08857_));
 AOI21_X2 _32556_ (.A(_08813_),
    .B1(_08825_),
    .B2(_08857_),
    .ZN(_08858_));
 XNOR2_X2 _32557_ (.A(_08827_),
    .B(_08858_),
    .ZN(_08859_));
 NAND2_X1 _32558_ (.A1(_08823_),
    .A2(_08814_),
    .ZN(_08860_));
 OAI21_X1 _32559_ (.A(_08835_),
    .B1(_08860_),
    .B2(_08839_),
    .ZN(_08861_));
 INV_X1 _32560_ (.A(_19990_),
    .ZN(_08862_));
 OAI21_X1 _32561_ (.A(_08756_),
    .B1(_08862_),
    .B2(_08758_),
    .ZN(_08863_));
 AOI21_X1 _32562_ (.A(_08755_),
    .B1(_08863_),
    .B2(_08760_),
    .ZN(_08864_));
 OAI21_X1 _32563_ (.A(_08754_),
    .B1(_08864_),
    .B2(_08762_),
    .ZN(_08865_));
 AOI21_X1 _32564_ (.A(_08753_),
    .B1(_08767_),
    .B2(_08865_),
    .ZN(_08866_));
 NOR3_X1 _32565_ (.A1(_08860_),
    .A2(_08840_),
    .A3(_08866_),
    .ZN(_08867_));
 OAI21_X1 _32566_ (.A(_08808_),
    .B1(_08861_),
    .B2(_08867_),
    .ZN(_08868_));
 NAND2_X1 _32567_ (.A1(_08833_),
    .A2(_08868_),
    .ZN(_08869_));
 AOI21_X1 _32568_ (.A(_19964_),
    .B1(_08869_),
    .B2(_08811_),
    .ZN(_08870_));
 OAI21_X1 _32569_ (.A(_08806_),
    .B1(_08807_),
    .B2(_08870_),
    .ZN(_08871_));
 AOI21_X1 _32570_ (.A(_19960_),
    .B1(_08871_),
    .B2(_08827_),
    .ZN(_08872_));
 XNOR2_X1 _32571_ (.A(_08804_),
    .B(_08872_),
    .ZN(_08873_));
 OR2_X1 _32572_ (.A1(_08816_),
    .A2(_08824_),
    .ZN(_08874_));
 OAI221_X1 _32573_ (.A(_08809_),
    .B1(_08815_),
    .B2(_08824_),
    .C1(_08874_),
    .C2(_08799_),
    .ZN(_08875_));
 XNOR2_X1 _32574_ (.A(_08822_),
    .B(_08875_),
    .ZN(_08876_));
 INV_X1 _32575_ (.A(_08876_),
    .ZN(_08877_));
 XNOR2_X1 _32576_ (.A(_08745_),
    .B(_08768_),
    .ZN(_08878_));
 AOI21_X1 _32577_ (.A(_08841_),
    .B1(_08842_),
    .B2(_08772_),
    .ZN(_08879_));
 XNOR2_X1 _32578_ (.A(_08814_),
    .B(_08879_),
    .ZN(_08880_));
 NAND3_X1 _32579_ (.A1(_08878_),
    .A2(_20007_),
    .A3(_08880_),
    .ZN(_08881_));
 NOR3_X1 _32580_ (.A1(_08768_),
    .A2(_08860_),
    .A3(_08840_),
    .ZN(_08882_));
 NOR2_X1 _32581_ (.A1(_08861_),
    .A2(_08882_),
    .ZN(_08883_));
 XNOR2_X1 _32582_ (.A(_08834_),
    .B(_08883_),
    .ZN(_08884_));
 XOR2_X2 _32583_ (.A(_08823_),
    .B(_08856_),
    .Z(_08885_));
 OR3_X1 _32584_ (.A1(_08881_),
    .A2(_08884_),
    .A3(_08885_),
    .ZN(_08886_));
 OAI21_X1 _32585_ (.A(_08837_),
    .B1(_08838_),
    .B2(_08879_),
    .ZN(_08887_));
 XNOR2_X2 _32586_ (.A(_19963_),
    .B(_08887_),
    .ZN(_08888_));
 NOR3_X1 _32587_ (.A1(_08877_),
    .A2(_08886_),
    .A3(_08888_),
    .ZN(_08889_));
 AND3_X1 _32588_ (.A1(_08859_),
    .A2(_08873_),
    .A3(_08889_),
    .ZN(_08890_));
 INV_X1 _32589_ (.A(_19958_),
    .ZN(_08891_));
 INV_X1 _32590_ (.A(_08804_),
    .ZN(_08892_));
 AOI21_X1 _32591_ (.A(_08755_),
    .B1(_19988_),
    .B2(_08760_),
    .ZN(_08893_));
 OAI21_X1 _32592_ (.A(_08796_),
    .B1(_08797_),
    .B2(_08893_),
    .ZN(_08894_));
 AOI21_X1 _32593_ (.A(_08794_),
    .B1(_08795_),
    .B2(_08894_),
    .ZN(_08895_));
 OAI221_X1 _32594_ (.A(_08809_),
    .B1(_08815_),
    .B2(_08824_),
    .C1(_08874_),
    .C2(_08895_),
    .ZN(_08896_));
 AOI21_X1 _32595_ (.A(_19964_),
    .B1(_08896_),
    .B2(_08811_),
    .ZN(_08897_));
 OAI21_X1 _32596_ (.A(_08806_),
    .B1(_08807_),
    .B2(_08897_),
    .ZN(_08898_));
 AOI21_X1 _32597_ (.A(_19960_),
    .B1(_08898_),
    .B2(_08827_),
    .ZN(_08899_));
 OAI21_X1 _32598_ (.A(_08891_),
    .B1(_08892_),
    .B2(_08899_),
    .ZN(_08900_));
 XNOR2_X2 _32599_ (.A(_08803_),
    .B(_08900_),
    .ZN(_08901_));
 NAND2_X1 _32600_ (.A1(_08890_),
    .A2(_08901_),
    .ZN(_08902_));
 NOR2_X1 _32601_ (.A1(_08853_),
    .A2(_08902_),
    .ZN(_08903_));
 XOR2_X1 _32602_ (.A(_08832_),
    .B(_08903_),
    .Z(_14382_));
 OR4_X1 _32603_ (.A1(\g_row[2].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08904_));
 OAI21_X2 _32604_ (.A(_07176_),
    .B1(_08904_),
    .B2(\g_row[2].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08905_));
 AND4_X1 _32605_ (.A1(\g_row[2].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_08906_));
 AOI21_X4 _32606_ (.A(_07180_),
    .B1(_08906_),
    .B2(\g_row[2].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_08907_));
 INV_X1 _32607_ (.A(_14380_),
    .ZN(_08908_));
 AOI21_X1 _32608_ (.A(_08905_),
    .B1(_08907_),
    .B2(_08908_),
    .ZN(_00337_));
 INV_X1 _32609_ (.A(_19997_),
    .ZN(_08909_));
 AOI21_X1 _32610_ (.A(_08905_),
    .B1(_08907_),
    .B2(_08909_),
    .ZN(_00338_));
 INV_X1 _32611_ (.A(_14388_),
    .ZN(_08910_));
 AOI21_X1 _32612_ (.A(_08905_),
    .B1(_08907_),
    .B2(_08910_),
    .ZN(_00339_));
 XOR2_X1 _32613_ (.A(_14387_),
    .B(_20006_),
    .Z(_08911_));
 AOI21_X1 _32614_ (.A(_08905_),
    .B1(_08907_),
    .B2(_08911_),
    .ZN(_00340_));
 AOI21_X1 _32615_ (.A(_20001_),
    .B1(_20002_),
    .B2(_19996_),
    .ZN(_08912_));
 INV_X1 _32616_ (.A(_08912_),
    .ZN(_08913_));
 AOI21_X1 _32617_ (.A(_20005_),
    .B1(_08913_),
    .B2(_20006_),
    .ZN(_08914_));
 XNOR2_X1 _32618_ (.A(\g_row[2].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20003_),
    .ZN(_08915_));
 XNOR2_X1 _32619_ (.A(_07174_),
    .B(_08915_),
    .ZN(_08916_));
 XNOR2_X1 _32620_ (.A(_08914_),
    .B(_08916_),
    .ZN(_08917_));
 AOI21_X1 _32621_ (.A(_08905_),
    .B1(_08907_),
    .B2(_08917_),
    .ZN(_00341_));
 INV_X1 _32622_ (.A(_08905_),
    .ZN(_08918_));
 NAND2_X4 _32623_ (.A1(_08918_),
    .A2(_08907_),
    .ZN(_08919_));
 INV_X1 _32624_ (.A(_14382_),
    .ZN(_14378_));
 NAND2_X1 _32625_ (.A1(_20010_),
    .A2(_14378_),
    .ZN(_08920_));
 NAND3_X1 _32626_ (.A1(_08878_),
    .A2(_08801_),
    .A3(_14382_),
    .ZN(_08921_));
 AOI21_X1 _32627_ (.A(_08919_),
    .B1(_08920_),
    .B2(_08921_),
    .ZN(_00336_));
 XNOR2_X1 _32628_ (.A(_20009_),
    .B(_08880_),
    .ZN(_08922_));
 INV_X1 _32629_ (.A(_20010_),
    .ZN(_08923_));
 MUX2_X1 _32630_ (.A(_08922_),
    .B(_08923_),
    .S(_14382_),
    .Z(_08924_));
 NOR2_X1 _32631_ (.A1(_08919_),
    .A2(_08924_),
    .ZN(_00342_));
 XNOR2_X1 _32632_ (.A(_08881_),
    .B(_08885_),
    .ZN(_08925_));
 MUX2_X1 _32633_ (.A(_08925_),
    .B(_08922_),
    .S(_14382_),
    .Z(_08926_));
 NOR2_X1 _32634_ (.A1(_08919_),
    .A2(_08926_),
    .ZN(_00343_));
 INV_X1 _32635_ (.A(_08884_),
    .ZN(_08927_));
 INV_X1 _32636_ (.A(_08885_),
    .ZN(_08928_));
 AND3_X1 _32637_ (.A1(_20009_),
    .A2(_08880_),
    .A3(_08928_),
    .ZN(_08929_));
 XNOR2_X1 _32638_ (.A(_08927_),
    .B(_08929_),
    .ZN(_08930_));
 MUX2_X1 _32639_ (.A(_08930_),
    .B(_08925_),
    .S(_14382_),
    .Z(_08931_));
 NOR2_X1 _32640_ (.A1(_08919_),
    .A2(_08931_),
    .ZN(_00344_));
 XNOR2_X1 _32641_ (.A(_08877_),
    .B(_08886_),
    .ZN(_08932_));
 MUX2_X1 _32642_ (.A(_08932_),
    .B(_08930_),
    .S(_14382_),
    .Z(_08933_));
 NOR2_X1 _32643_ (.A1(_08919_),
    .A2(_08933_),
    .ZN(_00345_));
 AND3_X1 _32644_ (.A1(_08876_),
    .A2(_08927_),
    .A3(_08929_),
    .ZN(_08934_));
 XOR2_X1 _32645_ (.A(_08888_),
    .B(_08934_),
    .Z(_08935_));
 MUX2_X1 _32646_ (.A(_08935_),
    .B(_08932_),
    .S(_14382_),
    .Z(_08936_));
 NOR2_X1 _32647_ (.A1(_08919_),
    .A2(_08936_),
    .ZN(_00346_));
 XNOR2_X1 _32648_ (.A(_08859_),
    .B(_08889_),
    .ZN(_08937_));
 MUX2_X1 _32649_ (.A(_08937_),
    .B(_08935_),
    .S(_14382_),
    .Z(_08938_));
 NOR2_X1 _32650_ (.A1(_08919_),
    .A2(_08938_),
    .ZN(_00347_));
 NAND2_X1 _32651_ (.A1(_08859_),
    .A2(_08934_),
    .ZN(_08939_));
 NOR2_X1 _32652_ (.A1(_08888_),
    .A2(_08939_),
    .ZN(_08940_));
 XNOR2_X1 _32653_ (.A(_08873_),
    .B(_08940_),
    .ZN(_08941_));
 MUX2_X1 _32654_ (.A(_08941_),
    .B(_08937_),
    .S(_14382_),
    .Z(_08942_));
 NOR2_X1 _32655_ (.A1(_08919_),
    .A2(_08942_),
    .ZN(_00348_));
 AND2_X1 _32656_ (.A1(_08890_),
    .A2(_08901_),
    .ZN(_08943_));
 AOI21_X1 _32657_ (.A(_08919_),
    .B1(_08941_),
    .B2(_08943_),
    .ZN(_08944_));
 NOR2_X1 _32658_ (.A1(_08890_),
    .A2(_08901_),
    .ZN(_08945_));
 AOI21_X1 _32659_ (.A(_08945_),
    .B1(_08943_),
    .B2(_08853_),
    .ZN(_08946_));
 OAI21_X1 _32660_ (.A(_08944_),
    .B1(_08946_),
    .B2(_08832_),
    .ZN(_08947_));
 OR2_X1 _32661_ (.A1(_08903_),
    .A2(_08941_),
    .ZN(_08948_));
 AOI21_X2 _32662_ (.A(_08947_),
    .B1(_08948_),
    .B2(_08832_),
    .ZN(_00349_));
 AND2_X1 _32663_ (.A1(_08873_),
    .A2(_08940_),
    .ZN(_08949_));
 OAI21_X1 _32664_ (.A(_08901_),
    .B1(_08949_),
    .B2(_08890_),
    .ZN(_08950_));
 NOR2_X1 _32665_ (.A1(_08853_),
    .A2(_08950_),
    .ZN(_08951_));
 NAND2_X1 _32666_ (.A1(_08901_),
    .A2(_08949_),
    .ZN(_08952_));
 AOI21_X1 _32667_ (.A(_08951_),
    .B1(_08952_),
    .B2(_08853_),
    .ZN(_08953_));
 OAI21_X1 _32668_ (.A(_08890_),
    .B1(_08853_),
    .B2(_08949_),
    .ZN(_08954_));
 MUX2_X1 _32669_ (.A(_08890_),
    .B(_08954_),
    .S(_08901_),
    .Z(_08955_));
 MUX2_X1 _32670_ (.A(_08953_),
    .B(_08955_),
    .S(_08832_),
    .Z(_08956_));
 AND3_X1 _32671_ (.A1(_08918_),
    .A2(_08907_),
    .A3(_08956_),
    .ZN(_00350_));
 CLKBUF_X2 _32672_ (.A(_20034_),
    .Z(_08957_));
 AOI21_X1 _32673_ (.A(_20033_),
    .B1(_08957_),
    .B2(_20035_),
    .ZN(_08958_));
 BUF_X1 _32674_ (.A(_20036_),
    .Z(_08959_));
 NAND2_X1 _32675_ (.A1(_08957_),
    .A2(_08959_),
    .ZN(_08960_));
 CLKBUF_X2 _32676_ (.A(_20039_),
    .Z(_08961_));
 AOI21_X1 _32677_ (.A(_20037_),
    .B1(_20038_),
    .B2(_08961_),
    .ZN(_08962_));
 OAI21_X1 _32678_ (.A(_08958_),
    .B1(_08960_),
    .B2(_08962_),
    .ZN(_08963_));
 INV_X1 _32679_ (.A(_20041_),
    .ZN(_08964_));
 CLKBUF_X2 _32680_ (.A(_20043_),
    .Z(_08965_));
 INV_X1 _32681_ (.A(_20045_),
    .ZN(_08966_));
 AOI21_X1 _32682_ (.A(_20047_),
    .B1(_20048_),
    .B2(_20049_),
    .ZN(_08967_));
 INV_X1 _32683_ (.A(_20046_),
    .ZN(_08968_));
 OAI21_X1 _32684_ (.A(_08966_),
    .B1(_08967_),
    .B2(_08968_),
    .ZN(_08969_));
 CLKBUF_X2 _32685_ (.A(_20044_),
    .Z(_08970_));
 AOI21_X1 _32686_ (.A(_08965_),
    .B1(_08969_),
    .B2(_08970_),
    .ZN(_08971_));
 INV_X1 _32687_ (.A(_20042_),
    .ZN(_08972_));
 OAI21_X2 _32688_ (.A(_08964_),
    .B1(_08971_),
    .B2(_08972_),
    .ZN(_08973_));
 INV_X1 _32689_ (.A(_20038_),
    .ZN(_08974_));
 CLKBUF_X2 _32690_ (.A(_20040_),
    .Z(_08975_));
 INV_X1 _32691_ (.A(_08975_),
    .ZN(_08976_));
 NOR3_X2 _32692_ (.A1(_08974_),
    .A2(_08976_),
    .A3(_08960_),
    .ZN(_08977_));
 AOI21_X2 _32693_ (.A(_08963_),
    .B1(_08973_),
    .B2(_08977_),
    .ZN(_08978_));
 XNOR2_X2 _32694_ (.A(_20032_),
    .B(_08978_),
    .ZN(_08979_));
 INV_X1 _32695_ (.A(_08979_),
    .ZN(_08980_));
 INV_X1 _32696_ (.A(_20037_),
    .ZN(_08981_));
 AOI21_X1 _32697_ (.A(_08961_),
    .B1(_08975_),
    .B2(_08973_),
    .ZN(_08982_));
 OAI21_X2 _32698_ (.A(_08981_),
    .B1(_08982_),
    .B2(_08974_),
    .ZN(_08983_));
 XNOR2_X1 _32699_ (.A(_08959_),
    .B(_08983_),
    .ZN(_08984_));
 XNOR2_X1 _32700_ (.A(_08976_),
    .B(_08973_),
    .ZN(_08985_));
 INV_X1 _32701_ (.A(_20031_),
    .ZN(_08986_));
 INV_X1 _32702_ (.A(_20032_),
    .ZN(_08987_));
 AOI21_X1 _32703_ (.A(_20035_),
    .B1(_08959_),
    .B2(_20037_),
    .ZN(_08988_));
 INV_X1 _32704_ (.A(_08988_),
    .ZN(_08989_));
 AOI21_X1 _32705_ (.A(_20033_),
    .B1(_08989_),
    .B2(_08957_),
    .ZN(_08990_));
 OAI21_X1 _32706_ (.A(_08986_),
    .B1(_08987_),
    .B2(_08990_),
    .ZN(_08991_));
 INV_X1 _32707_ (.A(_08957_),
    .ZN(_08992_));
 NAND2_X1 _32708_ (.A1(_08959_),
    .A2(_20038_),
    .ZN(_08993_));
 NOR3_X2 _32709_ (.A1(_08987_),
    .A2(_08992_),
    .A3(_08993_),
    .ZN(_08994_));
 AOI21_X2 _32710_ (.A(_08961_),
    .B1(_08975_),
    .B2(_20041_),
    .ZN(_08995_));
 OAI21_X1 _32711_ (.A(_08966_),
    .B1(_08968_),
    .B2(_14392_),
    .ZN(_08996_));
 AOI21_X1 _32712_ (.A(_08965_),
    .B1(_08996_),
    .B2(_08970_),
    .ZN(_08997_));
 NAND2_X1 _32713_ (.A1(_08975_),
    .A2(_20042_),
    .ZN(_08998_));
 NOR2_X1 _32714_ (.A1(_08997_),
    .A2(_08998_),
    .ZN(_08999_));
 INV_X1 _32715_ (.A(_08999_),
    .ZN(_09000_));
 NAND2_X1 _32716_ (.A1(_08995_),
    .A2(_09000_),
    .ZN(_09001_));
 AOI21_X1 _32717_ (.A(_08991_),
    .B1(_08994_),
    .B2(_09001_),
    .ZN(_09002_));
 XNOR2_X1 _32718_ (.A(_20030_),
    .B(_09002_),
    .ZN(_20064_));
 AOI21_X1 _32719_ (.A(_08976_),
    .B1(_08972_),
    .B2(_08964_),
    .ZN(_09003_));
 NOR2_X1 _32720_ (.A1(_08961_),
    .A2(_09003_),
    .ZN(_09004_));
 XNOR2_X1 _32721_ (.A(_08974_),
    .B(_09004_),
    .ZN(_09005_));
 XNOR2_X1 _32722_ (.A(_14392_),
    .B(_20046_),
    .ZN(_09006_));
 NOR4_X1 _32723_ (.A1(_14393_),
    .A2(\g_row[2].g_col[2].mult.adder.a[0] ),
    .A3(_20050_),
    .A4(_09006_),
    .ZN(_09007_));
 XNOR2_X1 _32724_ (.A(_08972_),
    .B(_08997_),
    .ZN(_09008_));
 XNOR2_X1 _32725_ (.A(_08970_),
    .B(_08969_),
    .ZN(_09009_));
 NAND4_X1 _32726_ (.A1(_09005_),
    .A2(_09007_),
    .A3(_09008_),
    .A4(_09009_),
    .ZN(_09010_));
 OAI21_X1 _32727_ (.A(_08988_),
    .B1(_08993_),
    .B2(_08995_),
    .ZN(_09011_));
 NOR2_X1 _32728_ (.A1(_08993_),
    .A2(_09000_),
    .ZN(_09012_));
 NOR2_X1 _32729_ (.A1(_09011_),
    .A2(_09012_),
    .ZN(_09013_));
 XNOR2_X1 _32730_ (.A(_08957_),
    .B(_09013_),
    .ZN(_09014_));
 NOR4_X1 _32731_ (.A1(_08985_),
    .A2(_20064_),
    .A3(_09010_),
    .A4(_09014_),
    .ZN(_09015_));
 AND2_X1 _32732_ (.A1(_08984_),
    .A2(_09015_),
    .ZN(_09016_));
 NOR2_X1 _32733_ (.A1(_08980_),
    .A2(_09016_),
    .ZN(_20065_));
 INV_X1 _32734_ (.A(_20011_),
    .ZN(_09017_));
 INV_X1 _32735_ (.A(_20012_),
    .ZN(_09018_));
 BUF_X2 _32736_ (.A(_20014_),
    .Z(_09019_));
 INV_X1 _32737_ (.A(_20015_),
    .ZN(_09020_));
 INV_X1 _32738_ (.A(_20016_),
    .ZN(_09021_));
 INV_X1 _32739_ (.A(_20021_),
    .ZN(_09022_));
 BUF_X2 _32740_ (.A(_20024_),
    .Z(_09023_));
 AOI21_X2 _32741_ (.A(_20023_),
    .B1(_09023_),
    .B2(_20025_),
    .ZN(_09024_));
 CLKBUF_X2 _32742_ (.A(_20022_),
    .Z(_09025_));
 INV_X1 _32743_ (.A(_09025_),
    .ZN(_09026_));
 OAI21_X1 _32744_ (.A(_09022_),
    .B1(_09024_),
    .B2(_09026_),
    .ZN(_09027_));
 AOI21_X1 _32745_ (.A(_20019_),
    .B1(_20020_),
    .B2(_09027_),
    .ZN(_09028_));
 BUF_X2 _32746_ (.A(_20028_),
    .Z(_09029_));
 AND2_X1 _32747_ (.A1(_09029_),
    .A2(_20030_),
    .ZN(_09030_));
 AOI21_X1 _32748_ (.A(_20033_),
    .B1(_09011_),
    .B2(_08957_),
    .ZN(_09031_));
 OAI21_X1 _32749_ (.A(_08986_),
    .B1(_08987_),
    .B2(_09031_),
    .ZN(_09032_));
 AOI221_X2 _32750_ (.A(_20027_),
    .B1(_09029_),
    .B2(_20029_),
    .C1(_09030_),
    .C2(_09032_),
    .ZN(_09033_));
 BUF_X2 _32751_ (.A(_20026_),
    .Z(_09034_));
 NAND4_X1 _32752_ (.A1(_20020_),
    .A2(_09025_),
    .A3(_09023_),
    .A4(_09034_),
    .ZN(_09035_));
 OAI21_X1 _32753_ (.A(_09028_),
    .B1(_09033_),
    .B2(_09035_),
    .ZN(_09036_));
 BUF_X2 _32754_ (.A(_20018_),
    .Z(_09037_));
 AOI21_X1 _32755_ (.A(_20017_),
    .B1(_09036_),
    .B2(_09037_),
    .ZN(_09038_));
 OAI21_X1 _32756_ (.A(_09020_),
    .B1(_09021_),
    .B2(_09038_),
    .ZN(_09039_));
 AOI21_X2 _32757_ (.A(_20013_),
    .B1(_09019_),
    .B2(_09039_),
    .ZN(_09040_));
 OAI21_X4 _32758_ (.A(_09017_),
    .B1(_09018_),
    .B2(_09040_),
    .ZN(_09041_));
 INV_X1 _32759_ (.A(_20023_),
    .ZN(_09042_));
 INV_X1 _32760_ (.A(_09023_),
    .ZN(_09043_));
 AOI21_X1 _32761_ (.A(_20025_),
    .B1(_09034_),
    .B2(_20027_),
    .ZN(_09044_));
 OAI21_X1 _32762_ (.A(_09042_),
    .B1(_09043_),
    .B2(_09044_),
    .ZN(_09045_));
 AOI21_X1 _32763_ (.A(_20021_),
    .B1(_09045_),
    .B2(_09025_),
    .ZN(_09046_));
 NAND4_X1 _32764_ (.A1(_09025_),
    .A2(_09023_),
    .A3(_09034_),
    .A4(_09029_),
    .ZN(_09047_));
 AOI21_X1 _32765_ (.A(_20029_),
    .B1(_20030_),
    .B2(_20031_),
    .ZN(_09048_));
 NAND2_X1 _32766_ (.A1(_20030_),
    .A2(_20032_),
    .ZN(_09049_));
 OAI21_X1 _32767_ (.A(_09048_),
    .B1(_09049_),
    .B2(_08958_),
    .ZN(_09050_));
 NOR2_X1 _32768_ (.A1(_08960_),
    .A2(_09049_),
    .ZN(_09051_));
 INV_X1 _32769_ (.A(_08965_),
    .ZN(_09052_));
 OAI21_X1 _32770_ (.A(_08964_),
    .B1(_09052_),
    .B2(_08972_),
    .ZN(_09053_));
 AOI21_X1 _32771_ (.A(_08961_),
    .B1(_08975_),
    .B2(_09053_),
    .ZN(_09054_));
 OAI21_X1 _32772_ (.A(_08981_),
    .B1(_09054_),
    .B2(_08974_),
    .ZN(_09055_));
 AOI21_X1 _32773_ (.A(_09050_),
    .B1(_09051_),
    .B2(_09055_),
    .ZN(_09056_));
 OAI21_X1 _32774_ (.A(_09046_),
    .B1(_09047_),
    .B2(_09056_),
    .ZN(_09057_));
 AOI21_X1 _32775_ (.A(_20019_),
    .B1(_20020_),
    .B2(_09057_),
    .ZN(_09058_));
 INV_X1 _32776_ (.A(_09058_),
    .ZN(_09059_));
 AOI21_X1 _32777_ (.A(_20017_),
    .B1(_09059_),
    .B2(_09037_),
    .ZN(_09060_));
 OAI21_X1 _32778_ (.A(_09020_),
    .B1(_09021_),
    .B2(_09060_),
    .ZN(_09061_));
 AOI21_X1 _32779_ (.A(_20013_),
    .B1(_09019_),
    .B2(_09061_),
    .ZN(_09062_));
 XNOR2_X1 _32780_ (.A(_20012_),
    .B(_09062_),
    .ZN(_09063_));
 INV_X1 _32781_ (.A(_09063_),
    .ZN(_09064_));
 INV_X1 _32782_ (.A(_20019_),
    .ZN(_09065_));
 INV_X1 _32783_ (.A(_20020_),
    .ZN(_09066_));
 AOI21_X2 _32784_ (.A(_20027_),
    .B1(_09029_),
    .B2(_20029_),
    .ZN(_09067_));
 NAND2_X1 _32785_ (.A1(_09023_),
    .A2(_09034_),
    .ZN(_09068_));
 NAND3_X1 _32786_ (.A1(_09023_),
    .A2(_09034_),
    .A3(_09030_),
    .ZN(_09069_));
 AOI21_X1 _32787_ (.A(_08965_),
    .B1(_20045_),
    .B2(_08970_),
    .ZN(_09070_));
 OAI21_X1 _32788_ (.A(_08995_),
    .B1(_08998_),
    .B2(_09070_),
    .ZN(_09071_));
 AOI21_X1 _32789_ (.A(_08991_),
    .B1(_08994_),
    .B2(_09071_),
    .ZN(_09072_));
 OAI221_X1 _32790_ (.A(_09024_),
    .B1(_09067_),
    .B2(_09068_),
    .C1(_09069_),
    .C2(_09072_),
    .ZN(_09073_));
 AOI21_X1 _32791_ (.A(_20021_),
    .B1(_09073_),
    .B2(_09025_),
    .ZN(_09074_));
 OAI21_X1 _32792_ (.A(_09065_),
    .B1(_09066_),
    .B2(_09074_),
    .ZN(_09075_));
 AOI21_X1 _32793_ (.A(_20017_),
    .B1(_09075_),
    .B2(_09037_),
    .ZN(_09076_));
 OAI21_X2 _32794_ (.A(_09020_),
    .B1(_09021_),
    .B2(_09076_),
    .ZN(_09077_));
 XNOR2_X2 _32795_ (.A(_09019_),
    .B(_09077_),
    .ZN(_09078_));
 NAND2_X1 _32796_ (.A1(_08994_),
    .A2(_09030_),
    .ZN(_09079_));
 OAI21_X2 _32797_ (.A(_09033_),
    .B1(_09079_),
    .B2(_09000_),
    .ZN(_09080_));
 INV_X1 _32798_ (.A(_09080_),
    .ZN(_09081_));
 OAI21_X1 _32799_ (.A(_09028_),
    .B1(_09035_),
    .B2(_09081_),
    .ZN(_09082_));
 XOR2_X2 _32800_ (.A(_09037_),
    .B(_09082_),
    .Z(_09083_));
 NAND2_X1 _32801_ (.A1(_09034_),
    .A2(_09029_),
    .ZN(_09084_));
 OAI21_X1 _32802_ (.A(_09044_),
    .B1(_09084_),
    .B2(_09048_),
    .ZN(_09085_));
 INV_X1 _32803_ (.A(_20047_),
    .ZN(_09086_));
 OAI21_X1 _32804_ (.A(_08966_),
    .B1(_09086_),
    .B2(_08968_),
    .ZN(_09087_));
 AOI21_X1 _32805_ (.A(_08965_),
    .B1(_09087_),
    .B2(_08970_),
    .ZN(_09088_));
 OAI21_X1 _32806_ (.A(_08964_),
    .B1(_09088_),
    .B2(_08972_),
    .ZN(_09089_));
 AOI21_X1 _32807_ (.A(_08963_),
    .B1(_08977_),
    .B2(_09089_),
    .ZN(_09090_));
 NOR3_X1 _32808_ (.A1(_09084_),
    .A2(_09049_),
    .A3(_09090_),
    .ZN(_09091_));
 OAI21_X1 _32809_ (.A(_09023_),
    .B1(_09085_),
    .B2(_09091_),
    .ZN(_09092_));
 NAND2_X1 _32810_ (.A1(_09042_),
    .A2(_09092_),
    .ZN(_09093_));
 AOI21_X1 _32811_ (.A(_20021_),
    .B1(_09093_),
    .B2(_09025_),
    .ZN(_09094_));
 OAI21_X1 _32812_ (.A(_09065_),
    .B1(_09066_),
    .B2(_09094_),
    .ZN(_09095_));
 AOI21_X2 _32813_ (.A(_20017_),
    .B1(_09095_),
    .B2(_09037_),
    .ZN(_09096_));
 XNOR2_X2 _32814_ (.A(_20016_),
    .B(_09096_),
    .ZN(_09097_));
 OAI221_X2 _32815_ (.A(_09024_),
    .B1(_09067_),
    .B2(_09068_),
    .C1(_09069_),
    .C2(_09002_),
    .ZN(_09098_));
 XNOR2_X2 _32816_ (.A(_09026_),
    .B(_09098_),
    .ZN(_09099_));
 AOI21_X2 _32817_ (.A(_09050_),
    .B1(_09051_),
    .B2(_08983_),
    .ZN(_09100_));
 XNOR2_X2 _32818_ (.A(_09029_),
    .B(_09100_),
    .ZN(_09101_));
 AND3_X1 _32819_ (.A1(_08979_),
    .A2(_20064_),
    .A3(_09101_),
    .ZN(_09102_));
 NOR3_X1 _32820_ (.A1(_08978_),
    .A2(_09084_),
    .A3(_09049_),
    .ZN(_09103_));
 NOR2_X1 _32821_ (.A1(_09085_),
    .A2(_09103_),
    .ZN(_09104_));
 XNOR2_X2 _32822_ (.A(_09043_),
    .B(_09104_),
    .ZN(_09105_));
 INV_X1 _32823_ (.A(_09105_),
    .ZN(_09106_));
 XOR2_X2 _32824_ (.A(_09034_),
    .B(_09080_),
    .Z(_09107_));
 AND3_X1 _32825_ (.A1(_09102_),
    .A2(_09106_),
    .A3(_09107_),
    .ZN(_09108_));
 OAI21_X1 _32826_ (.A(_09046_),
    .B1(_09047_),
    .B2(_09100_),
    .ZN(_09109_));
 XNOR2_X2 _32827_ (.A(_09066_),
    .B(_09109_),
    .ZN(_09110_));
 NAND3_X1 _32828_ (.A1(_09099_),
    .A2(_09108_),
    .A3(_09110_),
    .ZN(_09111_));
 INV_X1 _32829_ (.A(_09111_),
    .ZN(_09112_));
 NAND3_X1 _32830_ (.A1(_09083_),
    .A2(_09097_),
    .A3(_09112_),
    .ZN(_09113_));
 NOR3_X1 _32831_ (.A1(_09064_),
    .A2(_09078_),
    .A3(_09113_),
    .ZN(_09114_));
 XOR2_X1 _32832_ (.A(_09041_),
    .B(_09114_),
    .Z(_14395_));
 INV_X1 _32833_ (.A(_14395_),
    .ZN(_14398_));
 OR4_X2 _32834_ (.A1(\g_row[2].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09115_));
 OAI21_X4 _32835_ (.A(_07394_),
    .B1(_09115_),
    .B2(\g_row[2].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09116_));
 AND4_X1 _32836_ (.A1(\g_row[2].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09117_));
 AOI21_X4 _32837_ (.A(_07398_),
    .B1(_09117_),
    .B2(\g_row[2].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09118_));
 INV_X1 _32838_ (.A(_14397_),
    .ZN(_09119_));
 AOI21_X1 _32839_ (.A(_09116_),
    .B1(_09118_),
    .B2(_09119_),
    .ZN(_00353_));
 INV_X1 _32840_ (.A(_20054_),
    .ZN(_09120_));
 AOI21_X1 _32841_ (.A(_09116_),
    .B1(_09118_),
    .B2(_09120_),
    .ZN(_00354_));
 INV_X1 _32842_ (.A(_14405_),
    .ZN(_09121_));
 AOI21_X1 _32843_ (.A(_09116_),
    .B1(_09118_),
    .B2(_09121_),
    .ZN(_00355_));
 XOR2_X1 _32844_ (.A(_14404_),
    .B(_20063_),
    .Z(_09122_));
 AOI21_X1 _32845_ (.A(_09116_),
    .B1(_09118_),
    .B2(_09122_),
    .ZN(_00356_));
 AOI21_X1 _32846_ (.A(_20058_),
    .B1(_20059_),
    .B2(_20053_),
    .ZN(_09123_));
 INV_X1 _32847_ (.A(_09123_),
    .ZN(_09124_));
 AOI21_X1 _32848_ (.A(_20062_),
    .B1(_09124_),
    .B2(_20063_),
    .ZN(_09125_));
 XNOR2_X1 _32849_ (.A(\g_row[2].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20060_),
    .ZN(_09126_));
 XNOR2_X1 _32850_ (.A(_07392_),
    .B(_09126_),
    .ZN(_09127_));
 XNOR2_X1 _32851_ (.A(_09125_),
    .B(_09127_),
    .ZN(_09128_));
 AOI21_X1 _32852_ (.A(_09116_),
    .B1(_09118_),
    .B2(_09128_),
    .ZN(_00357_));
 INV_X1 _32853_ (.A(_09116_),
    .ZN(_09129_));
 NAND2_X4 _32854_ (.A1(_09129_),
    .A2(_09118_),
    .ZN(_09130_));
 NAND2_X1 _32855_ (.A1(_20067_),
    .A2(_14395_),
    .ZN(_09131_));
 NAND3_X1 _32856_ (.A1(_08979_),
    .A2(_09016_),
    .A3(_14398_),
    .ZN(_09132_));
 AOI21_X2 _32857_ (.A(_09130_),
    .B1(_09131_),
    .B2(_09132_),
    .ZN(_00352_));
 INV_X1 _32858_ (.A(_20067_),
    .ZN(_09133_));
 XNOR2_X1 _32859_ (.A(_20066_),
    .B(_09101_),
    .ZN(_09134_));
 MUX2_X1 _32860_ (.A(_09133_),
    .B(_09134_),
    .S(_14395_),
    .Z(_09135_));
 NOR2_X1 _32861_ (.A1(_09130_),
    .A2(_09135_),
    .ZN(_00358_));
 XNOR2_X1 _32862_ (.A(_09102_),
    .B(_09107_),
    .ZN(_09136_));
 MUX2_X1 _32863_ (.A(_09134_),
    .B(_09136_),
    .S(_14395_),
    .Z(_09137_));
 NOR2_X1 _32864_ (.A1(_09130_),
    .A2(_09137_),
    .ZN(_00359_));
 NAND3_X1 _32865_ (.A1(_20066_),
    .A2(_09101_),
    .A3(_09107_),
    .ZN(_09138_));
 XNOR2_X1 _32866_ (.A(_09105_),
    .B(_09138_),
    .ZN(_09139_));
 MUX2_X1 _32867_ (.A(_09136_),
    .B(_09139_),
    .S(_14395_),
    .Z(_09140_));
 NOR2_X1 _32868_ (.A1(_09130_),
    .A2(_09140_),
    .ZN(_00360_));
 XNOR2_X1 _32869_ (.A(_09099_),
    .B(_09108_),
    .ZN(_09141_));
 MUX2_X1 _32870_ (.A(_09139_),
    .B(_09141_),
    .S(_14395_),
    .Z(_09142_));
 NOR2_X1 _32871_ (.A1(_09130_),
    .A2(_09142_),
    .ZN(_00361_));
 INV_X1 _32872_ (.A(_09099_),
    .ZN(_09143_));
 NOR3_X1 _32873_ (.A1(_09143_),
    .A2(_09105_),
    .A3(_09138_),
    .ZN(_09144_));
 XNOR2_X1 _32874_ (.A(_09110_),
    .B(_09144_),
    .ZN(_09145_));
 MUX2_X1 _32875_ (.A(_09141_),
    .B(_09145_),
    .S(_14395_),
    .Z(_09146_));
 NOR2_X1 _32876_ (.A1(_09130_),
    .A2(_09146_),
    .ZN(_00362_));
 XOR2_X1 _32877_ (.A(_09083_),
    .B(_09111_),
    .Z(_09147_));
 MUX2_X1 _32878_ (.A(_09145_),
    .B(_09147_),
    .S(_14395_),
    .Z(_09148_));
 NOR2_X1 _32879_ (.A1(_09130_),
    .A2(_09148_),
    .ZN(_00363_));
 INV_X1 _32880_ (.A(_09097_),
    .ZN(_09149_));
 NAND3_X1 _32881_ (.A1(_09083_),
    .A2(_09110_),
    .A3(_09144_),
    .ZN(_09150_));
 XNOR2_X1 _32882_ (.A(_09149_),
    .B(_09150_),
    .ZN(_09151_));
 MUX2_X1 _32883_ (.A(_09147_),
    .B(_09151_),
    .S(_14395_),
    .Z(_09152_));
 NOR2_X1 _32884_ (.A1(_09130_),
    .A2(_09152_),
    .ZN(_00364_));
 AND3_X2 _32885_ (.A1(_09083_),
    .A2(_09097_),
    .A3(_09112_),
    .ZN(_09153_));
 XNOR2_X2 _32886_ (.A(_09153_),
    .B(_09078_),
    .ZN(_09154_));
 XOR2_X2 _32887_ (.A(_09019_),
    .B(_09077_),
    .Z(_09155_));
 NOR2_X1 _32888_ (.A1(_09153_),
    .A2(_09155_),
    .ZN(_09156_));
 NAND2_X1 _32889_ (.A1(_09041_),
    .A2(_09063_),
    .ZN(_09157_));
 OAI22_X2 _32890_ (.A1(_09041_),
    .A2(_09114_),
    .B1(_09156_),
    .B2(_09157_),
    .ZN(_09158_));
 INV_X1 _32891_ (.A(_09151_),
    .ZN(_09159_));
 AOI22_X4 _32892_ (.A1(_09041_),
    .A2(_09154_),
    .B1(_09158_),
    .B2(_09159_),
    .ZN(_09160_));
 NOR2_X1 _32893_ (.A1(_09130_),
    .A2(_09160_),
    .ZN(_00365_));
 NOR2_X1 _32894_ (.A1(_09149_),
    .A2(_09150_),
    .ZN(_09161_));
 NAND4_X1 _32895_ (.A1(_09041_),
    .A2(_09064_),
    .A3(_09155_),
    .A4(_09161_),
    .ZN(_09162_));
 OAI21_X1 _32896_ (.A(_09155_),
    .B1(_09161_),
    .B2(_09153_),
    .ZN(_09163_));
 NOR2_X1 _32897_ (.A1(_09041_),
    .A2(_09161_),
    .ZN(_09164_));
 AOI22_X2 _32898_ (.A1(_09041_),
    .A2(_09163_),
    .B1(_09164_),
    .B2(_09153_),
    .ZN(_09165_));
 XNOR2_X1 _32899_ (.A(_09153_),
    .B(_09155_),
    .ZN(_09166_));
 OAI221_X1 _32900_ (.A(_09162_),
    .B1(_09165_),
    .B2(_09064_),
    .C1(_09041_),
    .C2(_09166_),
    .ZN(_09167_));
 AND3_X1 _32901_ (.A1(_09129_),
    .A2(_09118_),
    .A3(_09167_),
    .ZN(_00366_));
 CLKBUF_X2 _32902_ (.A(_20091_),
    .Z(_09168_));
 AOI21_X1 _32903_ (.A(_20090_),
    .B1(_09168_),
    .B2(_20092_),
    .ZN(_09169_));
 BUF_X1 _32904_ (.A(_20093_),
    .Z(_09170_));
 NAND2_X1 _32905_ (.A1(_09168_),
    .A2(_09170_),
    .ZN(_09171_));
 CLKBUF_X2 _32906_ (.A(_20096_),
    .Z(_09172_));
 AOI21_X1 _32907_ (.A(_20094_),
    .B1(_20095_),
    .B2(_09172_),
    .ZN(_09173_));
 OAI21_X1 _32908_ (.A(_09169_),
    .B1(_09171_),
    .B2(_09173_),
    .ZN(_09174_));
 INV_X1 _32909_ (.A(_20098_),
    .ZN(_09175_));
 CLKBUF_X2 _32910_ (.A(_20100_),
    .Z(_09176_));
 INV_X1 _32911_ (.A(_20102_),
    .ZN(_09177_));
 AOI21_X1 _32912_ (.A(_20104_),
    .B1(_20105_),
    .B2(_20106_),
    .ZN(_09178_));
 INV_X1 _32913_ (.A(_20103_),
    .ZN(_09179_));
 OAI21_X1 _32914_ (.A(_09177_),
    .B1(_09178_),
    .B2(_09179_),
    .ZN(_09180_));
 CLKBUF_X2 _32915_ (.A(_20101_),
    .Z(_09181_));
 AOI21_X1 _32916_ (.A(_09176_),
    .B1(_09180_),
    .B2(_09181_),
    .ZN(_09182_));
 INV_X1 _32917_ (.A(_20099_),
    .ZN(_09183_));
 OAI21_X2 _32918_ (.A(_09175_),
    .B1(_09182_),
    .B2(_09183_),
    .ZN(_09184_));
 INV_X1 _32919_ (.A(_20095_),
    .ZN(_09185_));
 CLKBUF_X2 _32920_ (.A(_20097_),
    .Z(_09186_));
 INV_X1 _32921_ (.A(_09186_),
    .ZN(_09187_));
 NOR3_X2 _32922_ (.A1(_09185_),
    .A2(_09187_),
    .A3(_09171_),
    .ZN(_09188_));
 AOI21_X2 _32923_ (.A(_09174_),
    .B1(_09184_),
    .B2(_09188_),
    .ZN(_09189_));
 XNOR2_X2 _32924_ (.A(_20089_),
    .B(_09189_),
    .ZN(_09190_));
 INV_X1 _32925_ (.A(_09190_),
    .ZN(_09191_));
 INV_X1 _32926_ (.A(_20094_),
    .ZN(_09192_));
 AOI21_X1 _32927_ (.A(_09172_),
    .B1(_09186_),
    .B2(_09184_),
    .ZN(_09193_));
 OAI21_X2 _32928_ (.A(_09192_),
    .B1(_09193_),
    .B2(_09185_),
    .ZN(_09194_));
 XNOR2_X1 _32929_ (.A(_09170_),
    .B(_09194_),
    .ZN(_09195_));
 XNOR2_X1 _32930_ (.A(_09187_),
    .B(_09184_),
    .ZN(_09196_));
 INV_X1 _32931_ (.A(_20088_),
    .ZN(_09197_));
 INV_X1 _32932_ (.A(_20089_),
    .ZN(_09198_));
 AOI21_X1 _32933_ (.A(_20092_),
    .B1(_09170_),
    .B2(_20094_),
    .ZN(_09199_));
 INV_X1 _32934_ (.A(_09199_),
    .ZN(_09200_));
 AOI21_X1 _32935_ (.A(_20090_),
    .B1(_09200_),
    .B2(_09168_),
    .ZN(_09201_));
 OAI21_X1 _32936_ (.A(_09197_),
    .B1(_09198_),
    .B2(_09201_),
    .ZN(_09202_));
 INV_X1 _32937_ (.A(_09168_),
    .ZN(_09203_));
 NAND2_X1 _32938_ (.A1(_09170_),
    .A2(_20095_),
    .ZN(_09204_));
 NOR3_X2 _32939_ (.A1(_09198_),
    .A2(_09203_),
    .A3(_09204_),
    .ZN(_09205_));
 AOI21_X2 _32940_ (.A(_09172_),
    .B1(_09186_),
    .B2(_20098_),
    .ZN(_09206_));
 OAI21_X1 _32941_ (.A(_09177_),
    .B1(_09179_),
    .B2(_14409_),
    .ZN(_09207_));
 AOI21_X1 _32942_ (.A(_09176_),
    .B1(_09207_),
    .B2(_09181_),
    .ZN(_09208_));
 NAND2_X1 _32943_ (.A1(_09186_),
    .A2(_20099_),
    .ZN(_09209_));
 NOR2_X1 _32944_ (.A1(_09208_),
    .A2(_09209_),
    .ZN(_09210_));
 INV_X1 _32945_ (.A(_09210_),
    .ZN(_09211_));
 NAND2_X1 _32946_ (.A1(_09206_),
    .A2(_09211_),
    .ZN(_09212_));
 AOI21_X1 _32947_ (.A(_09202_),
    .B1(_09205_),
    .B2(_09212_),
    .ZN(_09213_));
 XNOR2_X1 _32948_ (.A(_20087_),
    .B(_09213_),
    .ZN(_20121_));
 AOI21_X1 _32949_ (.A(_09187_),
    .B1(_09183_),
    .B2(_09175_),
    .ZN(_09214_));
 NOR2_X1 _32950_ (.A1(_09172_),
    .A2(_09214_),
    .ZN(_09215_));
 XNOR2_X1 _32951_ (.A(_09185_),
    .B(_09215_),
    .ZN(_09216_));
 XNOR2_X1 _32952_ (.A(_14409_),
    .B(_20103_),
    .ZN(_09217_));
 NOR4_X1 _32953_ (.A1(_14410_),
    .A2(\g_row[2].g_col[3].mult.adder.a[0] ),
    .A3(_20107_),
    .A4(_09217_),
    .ZN(_09218_));
 XNOR2_X1 _32954_ (.A(_09183_),
    .B(_09208_),
    .ZN(_09219_));
 XNOR2_X1 _32955_ (.A(_09181_),
    .B(_09180_),
    .ZN(_09220_));
 NAND4_X1 _32956_ (.A1(_09216_),
    .A2(_09218_),
    .A3(_09219_),
    .A4(_09220_),
    .ZN(_09221_));
 OAI21_X1 _32957_ (.A(_09199_),
    .B1(_09204_),
    .B2(_09206_),
    .ZN(_09222_));
 NOR2_X1 _32958_ (.A1(_09204_),
    .A2(_09211_),
    .ZN(_09223_));
 NOR2_X1 _32959_ (.A1(_09222_),
    .A2(_09223_),
    .ZN(_09224_));
 XNOR2_X1 _32960_ (.A(_09168_),
    .B(_09224_),
    .ZN(_09225_));
 NOR4_X1 _32961_ (.A1(_09196_),
    .A2(_20121_),
    .A3(_09221_),
    .A4(_09225_),
    .ZN(_09226_));
 AND2_X1 _32962_ (.A1(_09195_),
    .A2(_09226_),
    .ZN(_09227_));
 NOR2_X1 _32963_ (.A1(_09191_),
    .A2(_09227_),
    .ZN(_20122_));
 INV_X1 _32964_ (.A(_20068_),
    .ZN(_09228_));
 INV_X1 _32965_ (.A(_20069_),
    .ZN(_09229_));
 BUF_X2 _32966_ (.A(_20071_),
    .Z(_09230_));
 INV_X1 _32967_ (.A(_20072_),
    .ZN(_09231_));
 INV_X1 _32968_ (.A(_20073_),
    .ZN(_09232_));
 INV_X1 _32969_ (.A(_20078_),
    .ZN(_09233_));
 BUF_X2 _32970_ (.A(_20081_),
    .Z(_09234_));
 AOI21_X2 _32971_ (.A(_20080_),
    .B1(_09234_),
    .B2(_20082_),
    .ZN(_09235_));
 CLKBUF_X2 _32972_ (.A(_20079_),
    .Z(_09236_));
 INV_X1 _32973_ (.A(_09236_),
    .ZN(_09237_));
 OAI21_X1 _32974_ (.A(_09233_),
    .B1(_09235_),
    .B2(_09237_),
    .ZN(_09238_));
 AOI21_X1 _32975_ (.A(_20076_),
    .B1(_20077_),
    .B2(_09238_),
    .ZN(_09239_));
 BUF_X2 _32976_ (.A(_20085_),
    .Z(_09240_));
 AND2_X1 _32977_ (.A1(_09240_),
    .A2(_20087_),
    .ZN(_09241_));
 AOI21_X1 _32978_ (.A(_20090_),
    .B1(_09222_),
    .B2(_09168_),
    .ZN(_09242_));
 OAI21_X1 _32979_ (.A(_09197_),
    .B1(_09198_),
    .B2(_09242_),
    .ZN(_09243_));
 AOI221_X2 _32980_ (.A(_20084_),
    .B1(_09240_),
    .B2(_20086_),
    .C1(_09241_),
    .C2(_09243_),
    .ZN(_09244_));
 BUF_X2 _32981_ (.A(_20083_),
    .Z(_09245_));
 NAND4_X1 _32982_ (.A1(_20077_),
    .A2(_09236_),
    .A3(_09234_),
    .A4(_09245_),
    .ZN(_09246_));
 OAI21_X1 _32983_ (.A(_09239_),
    .B1(_09244_),
    .B2(_09246_),
    .ZN(_09247_));
 BUF_X2 _32984_ (.A(_20075_),
    .Z(_09248_));
 AOI21_X1 _32985_ (.A(_20074_),
    .B1(_09247_),
    .B2(_09248_),
    .ZN(_09249_));
 OAI21_X1 _32986_ (.A(_09231_),
    .B1(_09232_),
    .B2(_09249_),
    .ZN(_09250_));
 AOI21_X2 _32987_ (.A(_20070_),
    .B1(_09230_),
    .B2(_09250_),
    .ZN(_09251_));
 OAI21_X4 _32988_ (.A(_09228_),
    .B1(_09229_),
    .B2(_09251_),
    .ZN(_09252_));
 INV_X1 _32989_ (.A(_20080_),
    .ZN(_09253_));
 INV_X1 _32990_ (.A(_09234_),
    .ZN(_09254_));
 AOI21_X1 _32991_ (.A(_20082_),
    .B1(_09245_),
    .B2(_20084_),
    .ZN(_09255_));
 OAI21_X1 _32992_ (.A(_09253_),
    .B1(_09254_),
    .B2(_09255_),
    .ZN(_09256_));
 AOI21_X1 _32993_ (.A(_20078_),
    .B1(_09256_),
    .B2(_09236_),
    .ZN(_09257_));
 NAND4_X1 _32994_ (.A1(_09236_),
    .A2(_09234_),
    .A3(_09245_),
    .A4(_09240_),
    .ZN(_09258_));
 AOI21_X1 _32995_ (.A(_20086_),
    .B1(_20087_),
    .B2(_20088_),
    .ZN(_09259_));
 NAND2_X1 _32996_ (.A1(_20087_),
    .A2(_20089_),
    .ZN(_09260_));
 OAI21_X1 _32997_ (.A(_09259_),
    .B1(_09260_),
    .B2(_09169_),
    .ZN(_09261_));
 NOR2_X1 _32998_ (.A1(_09171_),
    .A2(_09260_),
    .ZN(_09262_));
 INV_X1 _32999_ (.A(_09176_),
    .ZN(_09263_));
 OAI21_X1 _33000_ (.A(_09175_),
    .B1(_09263_),
    .B2(_09183_),
    .ZN(_09264_));
 AOI21_X1 _33001_ (.A(_09172_),
    .B1(_09186_),
    .B2(_09264_),
    .ZN(_09265_));
 OAI21_X1 _33002_ (.A(_09192_),
    .B1(_09265_),
    .B2(_09185_),
    .ZN(_09266_));
 AOI21_X1 _33003_ (.A(_09261_),
    .B1(_09262_),
    .B2(_09266_),
    .ZN(_09267_));
 OAI21_X1 _33004_ (.A(_09257_),
    .B1(_09258_),
    .B2(_09267_),
    .ZN(_09268_));
 AOI21_X1 _33005_ (.A(_20076_),
    .B1(_20077_),
    .B2(_09268_),
    .ZN(_09269_));
 INV_X1 _33006_ (.A(_09269_),
    .ZN(_09270_));
 AOI21_X1 _33007_ (.A(_20074_),
    .B1(_09270_),
    .B2(_09248_),
    .ZN(_09271_));
 OAI21_X1 _33008_ (.A(_09231_),
    .B1(_09232_),
    .B2(_09271_),
    .ZN(_09272_));
 AOI21_X2 _33009_ (.A(_20070_),
    .B1(_09230_),
    .B2(_09272_),
    .ZN(_09273_));
 XNOR2_X1 _33010_ (.A(_20069_),
    .B(_09273_),
    .ZN(_09274_));
 INV_X1 _33011_ (.A(_09274_),
    .ZN(_09275_));
 INV_X1 _33012_ (.A(_20076_),
    .ZN(_09276_));
 INV_X1 _33013_ (.A(_20077_),
    .ZN(_09277_));
 AOI21_X2 _33014_ (.A(_20084_),
    .B1(_09240_),
    .B2(_20086_),
    .ZN(_09278_));
 NAND2_X1 _33015_ (.A1(_09234_),
    .A2(_09245_),
    .ZN(_09279_));
 NAND3_X1 _33016_ (.A1(_09234_),
    .A2(_09245_),
    .A3(_09241_),
    .ZN(_09280_));
 AOI21_X1 _33017_ (.A(_09176_),
    .B1(_20102_),
    .B2(_09181_),
    .ZN(_09281_));
 OAI21_X1 _33018_ (.A(_09206_),
    .B1(_09209_),
    .B2(_09281_),
    .ZN(_09282_));
 AOI21_X1 _33019_ (.A(_09202_),
    .B1(_09205_),
    .B2(_09282_),
    .ZN(_09283_));
 OAI221_X1 _33020_ (.A(_09235_),
    .B1(_09278_),
    .B2(_09279_),
    .C1(_09280_),
    .C2(_09283_),
    .ZN(_09284_));
 AOI21_X1 _33021_ (.A(_20078_),
    .B1(_09284_),
    .B2(_09236_),
    .ZN(_09285_));
 OAI21_X1 _33022_ (.A(_09276_),
    .B1(_09277_),
    .B2(_09285_),
    .ZN(_09286_));
 AOI21_X2 _33023_ (.A(_20074_),
    .B1(_09286_),
    .B2(_09248_),
    .ZN(_09287_));
 OAI21_X4 _33024_ (.A(_09231_),
    .B1(_09232_),
    .B2(_09287_),
    .ZN(_09288_));
 XNOR2_X2 _33025_ (.A(_09230_),
    .B(_09288_),
    .ZN(_09289_));
 NAND2_X1 _33026_ (.A1(_09205_),
    .A2(_09241_),
    .ZN(_09290_));
 OAI21_X2 _33027_ (.A(_09244_),
    .B1(_09290_),
    .B2(_09211_),
    .ZN(_09291_));
 INV_X1 _33028_ (.A(_09291_),
    .ZN(_09292_));
 OAI21_X1 _33029_ (.A(_09239_),
    .B1(_09246_),
    .B2(_09292_),
    .ZN(_09293_));
 XOR2_X2 _33030_ (.A(_09248_),
    .B(_09293_),
    .Z(_09294_));
 NAND2_X1 _33031_ (.A1(_09245_),
    .A2(_09240_),
    .ZN(_09295_));
 OAI21_X1 _33032_ (.A(_09255_),
    .B1(_09295_),
    .B2(_09259_),
    .ZN(_09296_));
 INV_X1 _33033_ (.A(_20104_),
    .ZN(_09297_));
 OAI21_X1 _33034_ (.A(_09177_),
    .B1(_09297_),
    .B2(_09179_),
    .ZN(_09298_));
 AOI21_X1 _33035_ (.A(_09176_),
    .B1(_09298_),
    .B2(_09181_),
    .ZN(_09299_));
 OAI21_X1 _33036_ (.A(_09175_),
    .B1(_09299_),
    .B2(_09183_),
    .ZN(_09300_));
 AOI21_X1 _33037_ (.A(_09174_),
    .B1(_09188_),
    .B2(_09300_),
    .ZN(_09301_));
 NOR3_X1 _33038_ (.A1(_09295_),
    .A2(_09260_),
    .A3(_09301_),
    .ZN(_09302_));
 OAI21_X1 _33039_ (.A(_09234_),
    .B1(_09296_),
    .B2(_09302_),
    .ZN(_09303_));
 NAND2_X1 _33040_ (.A1(_09253_),
    .A2(_09303_),
    .ZN(_09304_));
 AOI21_X1 _33041_ (.A(_20078_),
    .B1(_09304_),
    .B2(_09236_),
    .ZN(_09305_));
 OAI21_X1 _33042_ (.A(_09276_),
    .B1(_09277_),
    .B2(_09305_),
    .ZN(_09306_));
 AOI21_X2 _33043_ (.A(_20074_),
    .B1(_09306_),
    .B2(_09248_),
    .ZN(_09307_));
 XNOR2_X2 _33044_ (.A(_20073_),
    .B(_09307_),
    .ZN(_09308_));
 OAI221_X2 _33045_ (.A(_09235_),
    .B1(_09278_),
    .B2(_09279_),
    .C1(_09280_),
    .C2(_09213_),
    .ZN(_09309_));
 XNOR2_X2 _33046_ (.A(_09237_),
    .B(_09309_),
    .ZN(_09310_));
 AOI21_X2 _33047_ (.A(_09261_),
    .B1(_09262_),
    .B2(_09194_),
    .ZN(_09311_));
 XNOR2_X2 _33048_ (.A(_09240_),
    .B(_09311_),
    .ZN(_09312_));
 AND3_X1 _33049_ (.A1(_09190_),
    .A2(_20121_),
    .A3(_09312_),
    .ZN(_09313_));
 NOR3_X1 _33050_ (.A1(_09189_),
    .A2(_09295_),
    .A3(_09260_),
    .ZN(_09314_));
 NOR2_X1 _33051_ (.A1(_09296_),
    .A2(_09314_),
    .ZN(_09315_));
 XNOR2_X2 _33052_ (.A(_09254_),
    .B(_09315_),
    .ZN(_09316_));
 INV_X1 _33053_ (.A(_09316_),
    .ZN(_09317_));
 XOR2_X2 _33054_ (.A(_09245_),
    .B(_09291_),
    .Z(_09318_));
 AND3_X1 _33055_ (.A1(_09313_),
    .A2(_09317_),
    .A3(_09318_),
    .ZN(_09319_));
 OAI21_X1 _33056_ (.A(_09257_),
    .B1(_09258_),
    .B2(_09311_),
    .ZN(_09320_));
 XNOR2_X2 _33057_ (.A(_09277_),
    .B(_09320_),
    .ZN(_09321_));
 NAND3_X1 _33058_ (.A1(_09310_),
    .A2(_09319_),
    .A3(_09321_),
    .ZN(_09322_));
 INV_X1 _33059_ (.A(_09322_),
    .ZN(_09323_));
 NAND3_X1 _33060_ (.A1(_09294_),
    .A2(_09308_),
    .A3(_09323_),
    .ZN(_09324_));
 NOR3_X1 _33061_ (.A1(_09275_),
    .A2(_09289_),
    .A3(_09324_),
    .ZN(_09325_));
 XOR2_X1 _33062_ (.A(_09252_),
    .B(_09325_),
    .Z(_14412_));
 INV_X1 _33063_ (.A(_14412_),
    .ZN(_14416_));
 OR4_X1 _33064_ (.A1(\g_row[2].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09326_));
 OAI21_X4 _33065_ (.A(_07621_),
    .B1(_09326_),
    .B2(\g_row[2].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09327_));
 AND4_X1 _33066_ (.A1(\g_row[2].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[2].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[2].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[2].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09328_));
 AOI21_X4 _33067_ (.A(_07625_),
    .B1(_09328_),
    .B2(\g_row[2].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09329_));
 INV_X1 _33068_ (.A(_14414_),
    .ZN(_09330_));
 AOI21_X1 _33069_ (.A(_09327_),
    .B1(_09329_),
    .B2(_09330_),
    .ZN(_00369_));
 INV_X1 _33070_ (.A(_20111_),
    .ZN(_09331_));
 AOI21_X1 _33071_ (.A(_09327_),
    .B1(_09329_),
    .B2(_09331_),
    .ZN(_00370_));
 INV_X1 _33072_ (.A(_14422_),
    .ZN(_09332_));
 AOI21_X1 _33073_ (.A(_09327_),
    .B1(_09329_),
    .B2(_09332_),
    .ZN(_00371_));
 XOR2_X1 _33074_ (.A(_14421_),
    .B(_20120_),
    .Z(_09333_));
 AOI21_X1 _33075_ (.A(_09327_),
    .B1(_09329_),
    .B2(_09333_),
    .ZN(_00372_));
 AOI21_X1 _33076_ (.A(_20115_),
    .B1(_20116_),
    .B2(_20110_),
    .ZN(_09334_));
 INV_X1 _33077_ (.A(_09334_),
    .ZN(_09335_));
 AOI21_X1 _33078_ (.A(_20119_),
    .B1(_09335_),
    .B2(_20120_),
    .ZN(_09336_));
 XNOR2_X1 _33079_ (.A(\g_row[2].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20117_),
    .ZN(_09337_));
 XNOR2_X1 _33080_ (.A(_07619_),
    .B(_09337_),
    .ZN(_09338_));
 XNOR2_X1 _33081_ (.A(_09336_),
    .B(_09338_),
    .ZN(_09339_));
 AOI21_X1 _33082_ (.A(_09327_),
    .B1(_09329_),
    .B2(_09339_),
    .ZN(_00373_));
 INV_X1 _33083_ (.A(_09327_),
    .ZN(_09340_));
 NAND2_X4 _33084_ (.A1(_09340_),
    .A2(_09329_),
    .ZN(_09341_));
 NAND2_X1 _33085_ (.A1(_20124_),
    .A2(_14412_),
    .ZN(_09342_));
 NAND3_X1 _33086_ (.A1(_09190_),
    .A2(_09227_),
    .A3(_14416_),
    .ZN(_09343_));
 AOI21_X1 _33087_ (.A(_09341_),
    .B1(_09342_),
    .B2(_09343_),
    .ZN(_00368_));
 INV_X1 _33088_ (.A(_20124_),
    .ZN(_09344_));
 XNOR2_X1 _33089_ (.A(_20123_),
    .B(_09312_),
    .ZN(_09345_));
 MUX2_X1 _33090_ (.A(_09344_),
    .B(_09345_),
    .S(_14412_),
    .Z(_09346_));
 NOR2_X1 _33091_ (.A1(_09341_),
    .A2(_09346_),
    .ZN(_00374_));
 XNOR2_X1 _33092_ (.A(_09313_),
    .B(_09318_),
    .ZN(_09347_));
 MUX2_X1 _33093_ (.A(_09345_),
    .B(_09347_),
    .S(_14412_),
    .Z(_09348_));
 NOR2_X1 _33094_ (.A1(_09341_),
    .A2(_09348_),
    .ZN(_00375_));
 NAND3_X1 _33095_ (.A1(_20123_),
    .A2(_09312_),
    .A3(_09318_),
    .ZN(_09349_));
 XNOR2_X1 _33096_ (.A(_09316_),
    .B(_09349_),
    .ZN(_09350_));
 MUX2_X1 _33097_ (.A(_09347_),
    .B(_09350_),
    .S(_14412_),
    .Z(_09351_));
 NOR2_X1 _33098_ (.A1(_09341_),
    .A2(_09351_),
    .ZN(_00376_));
 XNOR2_X1 _33099_ (.A(_09310_),
    .B(_09319_),
    .ZN(_09352_));
 MUX2_X1 _33100_ (.A(_09350_),
    .B(_09352_),
    .S(_14412_),
    .Z(_09353_));
 NOR2_X1 _33101_ (.A1(_09341_),
    .A2(_09353_),
    .ZN(_00377_));
 INV_X1 _33102_ (.A(_09310_),
    .ZN(_09354_));
 NOR3_X1 _33103_ (.A1(_09354_),
    .A2(_09316_),
    .A3(_09349_),
    .ZN(_09355_));
 XNOR2_X1 _33104_ (.A(_09321_),
    .B(_09355_),
    .ZN(_09356_));
 MUX2_X1 _33105_ (.A(_09352_),
    .B(_09356_),
    .S(_14412_),
    .Z(_09357_));
 NOR2_X1 _33106_ (.A1(_09341_),
    .A2(_09357_),
    .ZN(_00378_));
 XOR2_X1 _33107_ (.A(_09294_),
    .B(_09322_),
    .Z(_09358_));
 MUX2_X1 _33108_ (.A(_09356_),
    .B(_09358_),
    .S(_14412_),
    .Z(_09359_));
 NOR2_X1 _33109_ (.A1(_09341_),
    .A2(_09359_),
    .ZN(_00379_));
 INV_X1 _33110_ (.A(_09308_),
    .ZN(_09360_));
 NAND3_X1 _33111_ (.A1(_09294_),
    .A2(_09321_),
    .A3(_09355_),
    .ZN(_09361_));
 XNOR2_X1 _33112_ (.A(_09360_),
    .B(_09361_),
    .ZN(_09362_));
 MUX2_X1 _33113_ (.A(_09358_),
    .B(_09362_),
    .S(_14412_),
    .Z(_09363_));
 NOR2_X1 _33114_ (.A1(_09341_),
    .A2(_09363_),
    .ZN(_00380_));
 AND3_X2 _33115_ (.A1(_09294_),
    .A2(_09308_),
    .A3(_09323_),
    .ZN(_09364_));
 XNOR2_X1 _33116_ (.A(_09364_),
    .B(_09289_),
    .ZN(_09365_));
 XOR2_X2 _33117_ (.A(_09230_),
    .B(_09288_),
    .Z(_09366_));
 NOR2_X1 _33118_ (.A1(_09364_),
    .A2(_09366_),
    .ZN(_09367_));
 NAND2_X1 _33119_ (.A1(_09252_),
    .A2(_09274_),
    .ZN(_09368_));
 OAI22_X1 _33120_ (.A1(_09252_),
    .A2(_09325_),
    .B1(_09367_),
    .B2(_09368_),
    .ZN(_09369_));
 INV_X1 _33121_ (.A(_09362_),
    .ZN(_09370_));
 AOI22_X1 _33122_ (.A1(_09252_),
    .A2(_09365_),
    .B1(_09369_),
    .B2(_09370_),
    .ZN(_09371_));
 NOR2_X1 _33123_ (.A1(_09341_),
    .A2(_09371_),
    .ZN(_00381_));
 NOR2_X1 _33124_ (.A1(_09360_),
    .A2(_09361_),
    .ZN(_09372_));
 NAND4_X1 _33125_ (.A1(_09252_),
    .A2(_09275_),
    .A3(_09366_),
    .A4(_09372_),
    .ZN(_09373_));
 OAI21_X1 _33126_ (.A(_09366_),
    .B1(_09372_),
    .B2(_09364_),
    .ZN(_09374_));
 NOR2_X1 _33127_ (.A1(_09252_),
    .A2(_09372_),
    .ZN(_09375_));
 AOI22_X1 _33128_ (.A1(_09252_),
    .A2(_09374_),
    .B1(_09375_),
    .B2(_09364_),
    .ZN(_09376_));
 XNOR2_X1 _33129_ (.A(_09364_),
    .B(_09366_),
    .ZN(_09377_));
 OAI221_X2 _33130_ (.A(_09373_),
    .B1(_09376_),
    .B2(_09275_),
    .C1(_09252_),
    .C2(_09377_),
    .ZN(_09378_));
 AND3_X1 _33131_ (.A1(_09340_),
    .A2(_09329_),
    .A3(_09378_),
    .ZN(_00382_));
 INV_X1 _33132_ (.A(_20146_),
    .ZN(_09379_));
 CLKBUF_X2 _33133_ (.A(_20148_),
    .Z(_09380_));
 AOI21_X1 _33134_ (.A(_20147_),
    .B1(_09380_),
    .B2(_20149_),
    .ZN(_09381_));
 BUF_X1 _33135_ (.A(_20150_),
    .Z(_09382_));
 NAND2_X1 _33136_ (.A1(_09380_),
    .A2(_09382_),
    .ZN(_09383_));
 CLKBUF_X2 _33137_ (.A(_20153_),
    .Z(_09384_));
 AOI21_X1 _33138_ (.A(_20151_),
    .B1(_20152_),
    .B2(_09384_),
    .ZN(_09385_));
 OAI21_X1 _33139_ (.A(_09381_),
    .B1(_09383_),
    .B2(_09385_),
    .ZN(_09386_));
 INV_X1 _33140_ (.A(_20155_),
    .ZN(_09387_));
 CLKBUF_X2 _33141_ (.A(_20157_),
    .Z(_09388_));
 INV_X1 _33142_ (.A(_20159_),
    .ZN(_09389_));
 AOI21_X1 _33143_ (.A(_20161_),
    .B1(_20162_),
    .B2(_20163_),
    .ZN(_09390_));
 INV_X1 _33144_ (.A(_20160_),
    .ZN(_09391_));
 OAI21_X1 _33145_ (.A(_09389_),
    .B1(_09390_),
    .B2(_09391_),
    .ZN(_09392_));
 CLKBUF_X2 _33146_ (.A(_20158_),
    .Z(_09393_));
 AOI21_X1 _33147_ (.A(_09388_),
    .B1(_09392_),
    .B2(_09393_),
    .ZN(_09394_));
 INV_X1 _33148_ (.A(_20156_),
    .ZN(_09395_));
 OAI21_X2 _33149_ (.A(_09387_),
    .B1(_09394_),
    .B2(_09395_),
    .ZN(_09396_));
 INV_X1 _33150_ (.A(_20152_),
    .ZN(_09397_));
 BUF_X2 _33151_ (.A(_20154_),
    .Z(_09398_));
 INV_X1 _33152_ (.A(_09398_),
    .ZN(_09399_));
 NOR3_X2 _33153_ (.A1(_09397_),
    .A2(_09399_),
    .A3(_09383_),
    .ZN(_09400_));
 AOI21_X2 _33154_ (.A(_09386_),
    .B1(_09396_),
    .B2(_09400_),
    .ZN(_09401_));
 XNOR2_X1 _33155_ (.A(_09379_),
    .B(_09401_),
    .ZN(_09402_));
 INV_X1 _33156_ (.A(_20151_),
    .ZN(_09403_));
 AOI21_X1 _33157_ (.A(_09384_),
    .B1(_09398_),
    .B2(_09396_),
    .ZN(_09404_));
 OAI21_X2 _33158_ (.A(_09403_),
    .B1(_09404_),
    .B2(_09397_),
    .ZN(_09405_));
 XNOR2_X1 _33159_ (.A(_09382_),
    .B(_09405_),
    .ZN(_09406_));
 XNOR2_X1 _33160_ (.A(_09398_),
    .B(_09396_),
    .ZN(_09407_));
 INV_X1 _33161_ (.A(_20145_),
    .ZN(_09408_));
 AOI21_X1 _33162_ (.A(_20149_),
    .B1(_09382_),
    .B2(_20151_),
    .ZN(_09409_));
 INV_X1 _33163_ (.A(_09409_),
    .ZN(_09410_));
 AOI21_X1 _33164_ (.A(_20147_),
    .B1(_09410_),
    .B2(_09380_),
    .ZN(_09411_));
 OAI21_X1 _33165_ (.A(_09408_),
    .B1(_09379_),
    .B2(_09411_),
    .ZN(_09412_));
 INV_X1 _33166_ (.A(_09380_),
    .ZN(_09413_));
 NAND2_X1 _33167_ (.A1(_09382_),
    .A2(_20152_),
    .ZN(_09414_));
 NOR3_X2 _33168_ (.A1(_09379_),
    .A2(_09413_),
    .A3(_09414_),
    .ZN(_09415_));
 AOI21_X2 _33169_ (.A(_09384_),
    .B1(_09398_),
    .B2(_20155_),
    .ZN(_09416_));
 OAI21_X1 _33170_ (.A(_09389_),
    .B1(_09391_),
    .B2(_14426_),
    .ZN(_09417_));
 AOI21_X1 _33171_ (.A(_09388_),
    .B1(_09417_),
    .B2(_09393_),
    .ZN(_09418_));
 NAND2_X1 _33172_ (.A1(_09398_),
    .A2(_20156_),
    .ZN(_09419_));
 NOR2_X1 _33173_ (.A1(_09418_),
    .A2(_09419_),
    .ZN(_09420_));
 INV_X1 _33174_ (.A(_09420_),
    .ZN(_09421_));
 NAND2_X1 _33175_ (.A1(_09416_),
    .A2(_09421_),
    .ZN(_09422_));
 AOI21_X1 _33176_ (.A(_09412_),
    .B1(_09415_),
    .B2(_09422_),
    .ZN(_09423_));
 XNOR2_X1 _33177_ (.A(_20144_),
    .B(_09423_),
    .ZN(_20178_));
 XNOR2_X1 _33178_ (.A(_09395_),
    .B(_09418_),
    .ZN(_09424_));
 XNOR2_X1 _33179_ (.A(_09393_),
    .B(_09392_),
    .ZN(_09425_));
 AOI21_X1 _33180_ (.A(_09399_),
    .B1(_09395_),
    .B2(_09387_),
    .ZN(_09426_));
 NOR2_X1 _33181_ (.A1(_09384_),
    .A2(_09426_),
    .ZN(_09427_));
 XNOR2_X1 _33182_ (.A(_09397_),
    .B(_09427_),
    .ZN(_09428_));
 XNOR2_X1 _33183_ (.A(_14426_),
    .B(_20160_),
    .ZN(_09429_));
 NOR4_X1 _33184_ (.A1(_14427_),
    .A2(\g_row[3].g_col[0].mult.adder.a[0] ),
    .A3(_20164_),
    .A4(_09429_),
    .ZN(_09430_));
 NAND4_X1 _33185_ (.A1(_09424_),
    .A2(_09425_),
    .A3(_09428_),
    .A4(_09430_),
    .ZN(_09431_));
 OAI21_X1 _33186_ (.A(_09409_),
    .B1(_09414_),
    .B2(_09416_),
    .ZN(_09432_));
 NOR2_X1 _33187_ (.A1(_09414_),
    .A2(_09421_),
    .ZN(_09433_));
 NOR2_X1 _33188_ (.A1(_09432_),
    .A2(_09433_),
    .ZN(_09434_));
 XNOR2_X1 _33189_ (.A(_09380_),
    .B(_09434_),
    .ZN(_09435_));
 NOR3_X1 _33190_ (.A1(_20178_),
    .A2(_09431_),
    .A3(_09435_),
    .ZN(_09436_));
 AND3_X1 _33191_ (.A1(_09406_),
    .A2(_09407_),
    .A3(_09436_),
    .ZN(_09437_));
 NOR2_X1 _33192_ (.A1(_09402_),
    .A2(_09437_),
    .ZN(_20179_));
 INV_X1 _33193_ (.A(_20125_),
    .ZN(_09438_));
 INV_X1 _33194_ (.A(_20126_),
    .ZN(_09439_));
 INV_X1 _33195_ (.A(_20129_),
    .ZN(_09440_));
 INV_X1 _33196_ (.A(_20130_),
    .ZN(_09441_));
 INV_X1 _33197_ (.A(_20135_),
    .ZN(_09442_));
 BUF_X2 _33198_ (.A(_20138_),
    .Z(_09443_));
 AOI21_X2 _33199_ (.A(_20137_),
    .B1(_09443_),
    .B2(_20139_),
    .ZN(_09444_));
 CLKBUF_X2 _33200_ (.A(_20136_),
    .Z(_09445_));
 INV_X1 _33201_ (.A(_09445_),
    .ZN(_09446_));
 OAI21_X1 _33202_ (.A(_09442_),
    .B1(_09444_),
    .B2(_09446_),
    .ZN(_09447_));
 AOI21_X1 _33203_ (.A(_20133_),
    .B1(_20134_),
    .B2(_09447_),
    .ZN(_09448_));
 BUF_X2 _33204_ (.A(_20142_),
    .Z(_09449_));
 AND2_X1 _33205_ (.A1(_09449_),
    .A2(_20144_),
    .ZN(_09450_));
 AOI21_X1 _33206_ (.A(_20147_),
    .B1(_09432_),
    .B2(_09380_),
    .ZN(_09451_));
 OAI21_X1 _33207_ (.A(_09408_),
    .B1(_09379_),
    .B2(_09451_),
    .ZN(_09452_));
 AOI221_X2 _33208_ (.A(_20141_),
    .B1(_09449_),
    .B2(_20143_),
    .C1(_09450_),
    .C2(_09452_),
    .ZN(_09453_));
 BUF_X2 _33209_ (.A(_20140_),
    .Z(_09454_));
 NAND4_X1 _33210_ (.A1(_20134_),
    .A2(_09445_),
    .A3(_09443_),
    .A4(_09454_),
    .ZN(_09455_));
 OAI21_X1 _33211_ (.A(_09448_),
    .B1(_09453_),
    .B2(_09455_),
    .ZN(_09456_));
 BUF_X2 _33212_ (.A(_20132_),
    .Z(_09457_));
 AOI21_X1 _33213_ (.A(_20131_),
    .B1(_09456_),
    .B2(_09457_),
    .ZN(_09458_));
 OAI21_X1 _33214_ (.A(_09440_),
    .B1(_09441_),
    .B2(_09458_),
    .ZN(_09459_));
 AOI21_X2 _33215_ (.A(_20127_),
    .B1(_20128_),
    .B2(_09459_),
    .ZN(_09460_));
 OAI21_X4 _33216_ (.A(_09438_),
    .B1(_09439_),
    .B2(_09460_),
    .ZN(_09461_));
 INV_X1 _33217_ (.A(_20137_),
    .ZN(_09462_));
 INV_X1 _33218_ (.A(_09443_),
    .ZN(_09463_));
 AOI21_X1 _33219_ (.A(_20139_),
    .B1(_09454_),
    .B2(_20141_),
    .ZN(_09464_));
 OAI21_X1 _33220_ (.A(_09462_),
    .B1(_09463_),
    .B2(_09464_),
    .ZN(_09465_));
 AOI21_X1 _33221_ (.A(_20135_),
    .B1(_09465_),
    .B2(_09445_),
    .ZN(_09466_));
 NAND4_X1 _33222_ (.A1(_09445_),
    .A2(_09443_),
    .A3(_09454_),
    .A4(_09449_),
    .ZN(_09467_));
 AOI21_X1 _33223_ (.A(_20143_),
    .B1(_20144_),
    .B2(_20145_),
    .ZN(_09468_));
 NAND2_X1 _33224_ (.A1(_20144_),
    .A2(_20146_),
    .ZN(_09469_));
 OAI21_X1 _33225_ (.A(_09468_),
    .B1(_09469_),
    .B2(_09381_),
    .ZN(_09470_));
 NOR2_X1 _33226_ (.A1(_09383_),
    .A2(_09469_),
    .ZN(_09471_));
 INV_X1 _33227_ (.A(_09388_),
    .ZN(_09472_));
 OAI21_X1 _33228_ (.A(_09387_),
    .B1(_09472_),
    .B2(_09395_),
    .ZN(_09473_));
 AOI21_X1 _33229_ (.A(_09384_),
    .B1(_09398_),
    .B2(_09473_),
    .ZN(_09474_));
 OAI21_X1 _33230_ (.A(_09403_),
    .B1(_09474_),
    .B2(_09397_),
    .ZN(_09475_));
 AOI21_X1 _33231_ (.A(_09470_),
    .B1(_09471_),
    .B2(_09475_),
    .ZN(_09476_));
 OAI21_X1 _33232_ (.A(_09466_),
    .B1(_09467_),
    .B2(_09476_),
    .ZN(_09477_));
 AOI21_X1 _33233_ (.A(_20133_),
    .B1(_20134_),
    .B2(_09477_),
    .ZN(_09478_));
 INV_X1 _33234_ (.A(_09478_),
    .ZN(_09479_));
 AOI21_X1 _33235_ (.A(_20131_),
    .B1(_09479_),
    .B2(_09457_),
    .ZN(_09480_));
 OAI21_X1 _33236_ (.A(_09440_),
    .B1(_09441_),
    .B2(_09480_),
    .ZN(_09481_));
 AOI21_X2 _33237_ (.A(_20127_),
    .B1(_20128_),
    .B2(_09481_),
    .ZN(_09482_));
 XNOR2_X2 _33238_ (.A(_20126_),
    .B(_09482_),
    .ZN(_09483_));
 INV_X1 _33239_ (.A(_09483_),
    .ZN(_09484_));
 INV_X1 _33240_ (.A(_20133_),
    .ZN(_09485_));
 INV_X1 _33241_ (.A(_20134_),
    .ZN(_09486_));
 AOI21_X2 _33242_ (.A(_20141_),
    .B1(_09449_),
    .B2(_20143_),
    .ZN(_09487_));
 NAND2_X1 _33243_ (.A1(_09443_),
    .A2(_09454_),
    .ZN(_09488_));
 NAND3_X1 _33244_ (.A1(_09443_),
    .A2(_09454_),
    .A3(_09450_),
    .ZN(_09489_));
 AOI21_X1 _33245_ (.A(_09388_),
    .B1(_20159_),
    .B2(_09393_),
    .ZN(_09490_));
 OAI21_X1 _33246_ (.A(_09416_),
    .B1(_09419_),
    .B2(_09490_),
    .ZN(_09491_));
 AOI21_X1 _33247_ (.A(_09412_),
    .B1(_09415_),
    .B2(_09491_),
    .ZN(_09492_));
 OAI221_X1 _33248_ (.A(_09444_),
    .B1(_09487_),
    .B2(_09488_),
    .C1(_09489_),
    .C2(_09492_),
    .ZN(_09493_));
 AOI21_X1 _33249_ (.A(_20135_),
    .B1(_09493_),
    .B2(_09445_),
    .ZN(_09494_));
 OAI21_X1 _33250_ (.A(_09485_),
    .B1(_09486_),
    .B2(_09494_),
    .ZN(_09495_));
 AOI21_X1 _33251_ (.A(_20131_),
    .B1(_09495_),
    .B2(_09457_),
    .ZN(_09496_));
 OAI21_X1 _33252_ (.A(_09440_),
    .B1(_09441_),
    .B2(_09496_),
    .ZN(_09497_));
 XNOR2_X2 _33253_ (.A(_20128_),
    .B(_09497_),
    .ZN(_09498_));
 NAND2_X1 _33254_ (.A1(_09415_),
    .A2(_09450_),
    .ZN(_09499_));
 OAI21_X2 _33255_ (.A(_09453_),
    .B1(_09499_),
    .B2(_09421_),
    .ZN(_09500_));
 INV_X1 _33256_ (.A(_09500_),
    .ZN(_09501_));
 OAI21_X1 _33257_ (.A(_09448_),
    .B1(_09455_),
    .B2(_09501_),
    .ZN(_09502_));
 XOR2_X2 _33258_ (.A(_09457_),
    .B(_09502_),
    .Z(_09503_));
 NAND2_X1 _33259_ (.A1(_09454_),
    .A2(_09449_),
    .ZN(_09504_));
 OAI21_X1 _33260_ (.A(_09464_),
    .B1(_09504_),
    .B2(_09468_),
    .ZN(_09505_));
 INV_X1 _33261_ (.A(_20161_),
    .ZN(_09506_));
 OAI21_X1 _33262_ (.A(_09389_),
    .B1(_09506_),
    .B2(_09391_),
    .ZN(_09507_));
 AOI21_X1 _33263_ (.A(_09388_),
    .B1(_09507_),
    .B2(_09393_),
    .ZN(_09508_));
 OAI21_X1 _33264_ (.A(_09387_),
    .B1(_09508_),
    .B2(_09395_),
    .ZN(_09509_));
 AOI21_X1 _33265_ (.A(_09386_),
    .B1(_09400_),
    .B2(_09509_),
    .ZN(_09510_));
 NOR3_X1 _33266_ (.A1(_09504_),
    .A2(_09469_),
    .A3(_09510_),
    .ZN(_09511_));
 OAI21_X1 _33267_ (.A(_09443_),
    .B1(_09505_),
    .B2(_09511_),
    .ZN(_09512_));
 NAND2_X1 _33268_ (.A1(_09462_),
    .A2(_09512_),
    .ZN(_09513_));
 AOI21_X1 _33269_ (.A(_20135_),
    .B1(_09513_),
    .B2(_09445_),
    .ZN(_09514_));
 OAI21_X1 _33270_ (.A(_09485_),
    .B1(_09486_),
    .B2(_09514_),
    .ZN(_09515_));
 AOI21_X2 _33271_ (.A(_20131_),
    .B1(_09515_),
    .B2(_09457_),
    .ZN(_09516_));
 XNOR2_X2 _33272_ (.A(_20130_),
    .B(_09516_),
    .ZN(_09517_));
 OAI221_X2 _33273_ (.A(_09444_),
    .B1(_09487_),
    .B2(_09488_),
    .C1(_09489_),
    .C2(_09423_),
    .ZN(_09518_));
 XNOR2_X2 _33274_ (.A(_09446_),
    .B(_09518_),
    .ZN(_09519_));
 INV_X1 _33275_ (.A(_09402_),
    .ZN(_09520_));
 AOI21_X2 _33276_ (.A(_09470_),
    .B1(_09471_),
    .B2(_09405_),
    .ZN(_09521_));
 XNOR2_X2 _33277_ (.A(_09449_),
    .B(_09521_),
    .ZN(_09522_));
 AND3_X1 _33278_ (.A1(_09520_),
    .A2(_20178_),
    .A3(_09522_),
    .ZN(_09523_));
 NOR3_X1 _33279_ (.A1(_09401_),
    .A2(_09504_),
    .A3(_09469_),
    .ZN(_09524_));
 NOR2_X1 _33280_ (.A1(_09505_),
    .A2(_09524_),
    .ZN(_09525_));
 XNOR2_X2 _33281_ (.A(_09463_),
    .B(_09525_),
    .ZN(_09526_));
 INV_X1 _33282_ (.A(_09526_),
    .ZN(_09527_));
 XOR2_X2 _33283_ (.A(_09454_),
    .B(_09500_),
    .Z(_09528_));
 AND3_X1 _33284_ (.A1(_09523_),
    .A2(_09527_),
    .A3(_09528_),
    .ZN(_09529_));
 OAI21_X1 _33285_ (.A(_09466_),
    .B1(_09467_),
    .B2(_09521_),
    .ZN(_09530_));
 XNOR2_X2 _33286_ (.A(_09486_),
    .B(_09530_),
    .ZN(_09531_));
 NAND3_X1 _33287_ (.A1(_09519_),
    .A2(_09529_),
    .A3(_09531_),
    .ZN(_09532_));
 INV_X1 _33288_ (.A(_09532_),
    .ZN(_09533_));
 NAND3_X1 _33289_ (.A1(_09503_),
    .A2(_09517_),
    .A3(_09533_),
    .ZN(_09534_));
 NOR3_X1 _33290_ (.A1(_09484_),
    .A2(_09498_),
    .A3(_09534_),
    .ZN(_09535_));
 XOR2_X2 _33291_ (.A(_09461_),
    .B(_09535_),
    .Z(_09536_));
 BUF_X1 _33292_ (.A(_09536_),
    .Z(_14429_));
 INV_X1 _33293_ (.A(_14429_),
    .ZN(_14433_));
 OR4_X2 _33294_ (.A1(\g_row[3].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09537_));
 OAI21_X4 _33295_ (.A(_06947_),
    .B1(_09537_),
    .B2(\g_row[3].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09538_));
 AND4_X1 _33296_ (.A1(\g_row[3].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09539_));
 AOI21_X4 _33297_ (.A(_06951_),
    .B1(_09539_),
    .B2(\g_row[3].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09540_));
 INV_X1 _33298_ (.A(_14431_),
    .ZN(_09541_));
 AOI21_X1 _33299_ (.A(_09538_),
    .B1(_09540_),
    .B2(_09541_),
    .ZN(_00385_));
 INV_X1 _33300_ (.A(_20168_),
    .ZN(_09542_));
 AOI21_X1 _33301_ (.A(_09538_),
    .B1(_09540_),
    .B2(_09542_),
    .ZN(_00386_));
 INV_X1 _33302_ (.A(_14439_),
    .ZN(_09543_));
 AOI21_X1 _33303_ (.A(_09538_),
    .B1(_09540_),
    .B2(_09543_),
    .ZN(_00387_));
 XOR2_X1 _33304_ (.A(_14438_),
    .B(_20177_),
    .Z(_09544_));
 AOI21_X1 _33305_ (.A(_09538_),
    .B1(_09540_),
    .B2(_09544_),
    .ZN(_00388_));
 AOI21_X1 _33306_ (.A(_20172_),
    .B1(_20173_),
    .B2(_20167_),
    .ZN(_09545_));
 INV_X1 _33307_ (.A(_09545_),
    .ZN(_09546_));
 AOI21_X1 _33308_ (.A(_20176_),
    .B1(_09546_),
    .B2(_20177_),
    .ZN(_09547_));
 XNOR2_X1 _33309_ (.A(\g_row[3].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20174_),
    .ZN(_09548_));
 XNOR2_X1 _33310_ (.A(_06945_),
    .B(_09548_),
    .ZN(_09549_));
 XNOR2_X1 _33311_ (.A(_09547_),
    .B(_09549_),
    .ZN(_09550_));
 AOI21_X1 _33312_ (.A(_09538_),
    .B1(_09540_),
    .B2(_09550_),
    .ZN(_00389_));
 INV_X1 _33313_ (.A(_09538_),
    .ZN(_09551_));
 AND2_X1 _33314_ (.A1(_09520_),
    .A2(_09437_),
    .ZN(_09552_));
 MUX2_X1 _33315_ (.A(_09552_),
    .B(_20181_),
    .S(_09536_),
    .Z(_09553_));
 AND3_X1 _33316_ (.A1(_09551_),
    .A2(_09540_),
    .A3(_09553_),
    .ZN(_00384_));
 NAND2_X4 _33317_ (.A1(_09551_),
    .A2(_09540_),
    .ZN(_09554_));
 NOR2_X1 _33318_ (.A1(_20181_),
    .A2(_14429_),
    .ZN(_09555_));
 XNOR2_X1 _33319_ (.A(_20180_),
    .B(_09522_),
    .ZN(_09556_));
 AND2_X1 _33320_ (.A1(_14429_),
    .A2(_09556_),
    .ZN(_09557_));
 NOR3_X1 _33321_ (.A1(_09554_),
    .A2(_09555_),
    .A3(_09557_),
    .ZN(_00390_));
 XNOR2_X1 _33322_ (.A(_09523_),
    .B(_09528_),
    .ZN(_09558_));
 MUX2_X1 _33323_ (.A(_09556_),
    .B(_09558_),
    .S(_14429_),
    .Z(_09559_));
 NOR2_X1 _33324_ (.A1(_09554_),
    .A2(_09559_),
    .ZN(_00391_));
 NAND3_X1 _33325_ (.A1(_20180_),
    .A2(_09522_),
    .A3(_09528_),
    .ZN(_09560_));
 XNOR2_X1 _33326_ (.A(_09526_),
    .B(_09560_),
    .ZN(_09561_));
 MUX2_X1 _33327_ (.A(_09558_),
    .B(_09561_),
    .S(_14429_),
    .Z(_09562_));
 NOR2_X1 _33328_ (.A1(_09554_),
    .A2(_09562_),
    .ZN(_00392_));
 XNOR2_X1 _33329_ (.A(_09519_),
    .B(_09529_),
    .ZN(_09563_));
 MUX2_X1 _33330_ (.A(_09561_),
    .B(_09563_),
    .S(_14429_),
    .Z(_09564_));
 NOR2_X1 _33331_ (.A1(_09554_),
    .A2(_09564_),
    .ZN(_00393_));
 INV_X1 _33332_ (.A(_09519_),
    .ZN(_09565_));
 NOR3_X1 _33333_ (.A1(_09565_),
    .A2(_09526_),
    .A3(_09560_),
    .ZN(_09566_));
 XNOR2_X1 _33334_ (.A(_09531_),
    .B(_09566_),
    .ZN(_09567_));
 MUX2_X1 _33335_ (.A(_09563_),
    .B(_09567_),
    .S(_14429_),
    .Z(_09568_));
 NOR2_X1 _33336_ (.A1(_09554_),
    .A2(_09568_),
    .ZN(_00394_));
 XOR2_X1 _33337_ (.A(_09503_),
    .B(_09532_),
    .Z(_09569_));
 MUX2_X1 _33338_ (.A(_09567_),
    .B(_09569_),
    .S(_09536_),
    .Z(_09570_));
 NOR2_X1 _33339_ (.A1(_09554_),
    .A2(_09570_),
    .ZN(_00395_));
 NAND3_X2 _33340_ (.A1(_09503_),
    .A2(_09531_),
    .A3(_09566_),
    .ZN(_09571_));
 XNOR2_X2 _33341_ (.A(_09517_),
    .B(_09571_),
    .ZN(_09572_));
 NAND2_X1 _33342_ (.A1(_14429_),
    .A2(_09572_),
    .ZN(_09573_));
 OR2_X1 _33343_ (.A1(_14429_),
    .A2(_09569_),
    .ZN(_09574_));
 AOI21_X1 _33344_ (.A(_09554_),
    .B1(_09573_),
    .B2(_09574_),
    .ZN(_00396_));
 AND3_X1 _33345_ (.A1(_09503_),
    .A2(_09517_),
    .A3(_09533_),
    .ZN(_09575_));
 XNOR2_X1 _33346_ (.A(_09575_),
    .B(_09498_),
    .ZN(_09576_));
 NAND2_X1 _33347_ (.A1(_09498_),
    .A2(_09534_),
    .ZN(_09577_));
 NAND3_X1 _33348_ (.A1(_09461_),
    .A2(_09483_),
    .A3(_09577_),
    .ZN(_09578_));
 OAI21_X1 _33349_ (.A(_09578_),
    .B1(_09535_),
    .B2(_09461_),
    .ZN(_09579_));
 AOI22_X2 _33350_ (.A1(_09461_),
    .A2(_09576_),
    .B1(_09579_),
    .B2(_09572_),
    .ZN(_09580_));
 NOR2_X1 _33351_ (.A1(_09554_),
    .A2(_09580_),
    .ZN(_00397_));
 INV_X1 _33352_ (.A(_09517_),
    .ZN(_09581_));
 NOR2_X1 _33353_ (.A1(_09581_),
    .A2(_09571_),
    .ZN(_09582_));
 OAI21_X1 _33354_ (.A(_09575_),
    .B1(_09484_),
    .B2(_09582_),
    .ZN(_09583_));
 OAI21_X1 _33355_ (.A(_09577_),
    .B1(_09583_),
    .B2(_09498_),
    .ZN(_09584_));
 NOR4_X1 _33356_ (.A1(_09581_),
    .A2(_09483_),
    .A3(_09498_),
    .A4(_09571_),
    .ZN(_09585_));
 INV_X1 _33357_ (.A(_09498_),
    .ZN(_09586_));
 OAI21_X1 _33358_ (.A(_09586_),
    .B1(_09582_),
    .B2(_09575_),
    .ZN(_09587_));
 AOI21_X1 _33359_ (.A(_09585_),
    .B1(_09587_),
    .B2(_09483_),
    .ZN(_09588_));
 MUX2_X1 _33360_ (.A(_09584_),
    .B(_09588_),
    .S(_09461_),
    .Z(_09589_));
 NOR2_X1 _33361_ (.A1(_09554_),
    .A2(_09589_),
    .ZN(_00398_));
 BUF_X1 _33362_ (.A(_20203_),
    .Z(_09590_));
 INV_X1 _33363_ (.A(_09590_),
    .ZN(_09591_));
 BUF_X1 _33364_ (.A(_20205_),
    .Z(_09592_));
 AOI21_X1 _33365_ (.A(_20204_),
    .B1(_09592_),
    .B2(_20206_),
    .ZN(_09593_));
 BUF_X2 _33366_ (.A(_20207_),
    .Z(_09594_));
 NAND2_X2 _33367_ (.A1(_09592_),
    .A2(_09594_),
    .ZN(_09595_));
 CLKBUF_X2 _33368_ (.A(_20210_),
    .Z(_09596_));
 AOI21_X1 _33369_ (.A(_20208_),
    .B1(_20209_),
    .B2(_09596_),
    .ZN(_09597_));
 OAI21_X1 _33370_ (.A(_09593_),
    .B1(_09595_),
    .B2(_09597_),
    .ZN(_09598_));
 INV_X1 _33371_ (.A(_20212_),
    .ZN(_09599_));
 CLKBUF_X2 _33372_ (.A(_20214_),
    .Z(_09600_));
 INV_X1 _33373_ (.A(_20216_),
    .ZN(_09601_));
 AOI21_X1 _33374_ (.A(_20218_),
    .B1(_20219_),
    .B2(_20220_),
    .ZN(_09602_));
 INV_X1 _33375_ (.A(_20217_),
    .ZN(_09603_));
 OAI21_X1 _33376_ (.A(_09601_),
    .B1(_09602_),
    .B2(_09603_),
    .ZN(_09604_));
 CLKBUF_X2 _33377_ (.A(_20215_),
    .Z(_09605_));
 AOI21_X1 _33378_ (.A(_09600_),
    .B1(_09604_),
    .B2(_09605_),
    .ZN(_09606_));
 INV_X1 _33379_ (.A(_20213_),
    .ZN(_09607_));
 OAI21_X1 _33380_ (.A(_09599_),
    .B1(_09606_),
    .B2(_09607_),
    .ZN(_09608_));
 INV_X2 _33381_ (.A(_20209_),
    .ZN(_09609_));
 CLKBUF_X2 _33382_ (.A(_20211_),
    .Z(_09610_));
 INV_X1 _33383_ (.A(_09610_),
    .ZN(_09611_));
 NOR3_X2 _33384_ (.A1(_09609_),
    .A2(_09611_),
    .A3(_09595_),
    .ZN(_09612_));
 AOI21_X2 _33385_ (.A(_09598_),
    .B1(_09608_),
    .B2(_09612_),
    .ZN(_09613_));
 XNOR2_X1 _33386_ (.A(_09591_),
    .B(_09613_),
    .ZN(_09614_));
 INV_X1 _33387_ (.A(_20208_),
    .ZN(_09615_));
 AOI21_X1 _33388_ (.A(_09596_),
    .B1(_09610_),
    .B2(_09608_),
    .ZN(_09616_));
 OAI21_X1 _33389_ (.A(_09615_),
    .B1(_09616_),
    .B2(_09609_),
    .ZN(_09617_));
 XOR2_X2 _33390_ (.A(_09594_),
    .B(_09617_),
    .Z(_09618_));
 NAND2_X1 _33391_ (.A1(_09609_),
    .A2(_09615_),
    .ZN(_09619_));
 AOI21_X1 _33392_ (.A(_20206_),
    .B1(_09594_),
    .B2(_09619_),
    .ZN(_09620_));
 XNOR2_X1 _33393_ (.A(_09592_),
    .B(_09620_),
    .ZN(_09621_));
 XNOR2_X1 _33394_ (.A(_14443_),
    .B(_20217_),
    .ZN(_09622_));
 OR4_X1 _33395_ (.A1(_14444_),
    .A2(\g_row[3].g_col[1].mult.adder.a[0] ),
    .A3(_20221_),
    .A4(_09622_),
    .ZN(_09623_));
 OAI21_X1 _33396_ (.A(_09601_),
    .B1(_09603_),
    .B2(_14443_),
    .ZN(_09624_));
 AOI21_X2 _33397_ (.A(_09600_),
    .B1(_09624_),
    .B2(_09605_),
    .ZN(_09625_));
 XNOR2_X1 _33398_ (.A(_20213_),
    .B(_09625_),
    .ZN(_09626_));
 NOR3_X1 _33399_ (.A1(_09621_),
    .A2(_09623_),
    .A3(_09626_),
    .ZN(_09627_));
 AOI21_X1 _33400_ (.A(_09611_),
    .B1(_09607_),
    .B2(_09599_),
    .ZN(_09628_));
 NOR2_X1 _33401_ (.A1(_09596_),
    .A2(_09628_),
    .ZN(_09629_));
 XNOR2_X1 _33402_ (.A(_09609_),
    .B(_09629_),
    .ZN(_09630_));
 XNOR2_X1 _33403_ (.A(_09605_),
    .B(_09604_),
    .ZN(_09631_));
 NAND3_X1 _33404_ (.A1(_09627_),
    .A2(_09630_),
    .A3(_09631_),
    .ZN(_09632_));
 CLKBUF_X2 _33405_ (.A(_20201_),
    .Z(_09633_));
 INV_X1 _33406_ (.A(_20204_),
    .ZN(_09634_));
 AOI21_X1 _33407_ (.A(_20206_),
    .B1(_09594_),
    .B2(_20208_),
    .ZN(_09635_));
 INV_X1 _33408_ (.A(_09592_),
    .ZN(_09636_));
 OAI21_X1 _33409_ (.A(_09634_),
    .B1(_09635_),
    .B2(_09636_),
    .ZN(_09637_));
 AND2_X1 _33410_ (.A1(_09590_),
    .A2(_09637_),
    .ZN(_09638_));
 OR2_X1 _33411_ (.A1(_20202_),
    .A2(_09638_),
    .ZN(_09639_));
 NOR3_X2 _33412_ (.A1(_09591_),
    .A2(_09609_),
    .A3(_09595_),
    .ZN(_09640_));
 AOI21_X2 _33413_ (.A(_09596_),
    .B1(_09610_),
    .B2(_20212_),
    .ZN(_09641_));
 NAND2_X1 _33414_ (.A1(_09610_),
    .A2(_20213_),
    .ZN(_09642_));
 OAI21_X1 _33415_ (.A(_09641_),
    .B1(_09642_),
    .B2(_09625_),
    .ZN(_09643_));
 AOI21_X2 _33416_ (.A(_09639_),
    .B1(_09640_),
    .B2(_09643_),
    .ZN(_09644_));
 XNOR2_X2 _33417_ (.A(_09633_),
    .B(_09644_),
    .ZN(_20235_));
 XNOR2_X1 _33418_ (.A(_09611_),
    .B(_09608_),
    .ZN(_09645_));
 NOR4_X1 _33419_ (.A1(_09618_),
    .A2(_09632_),
    .A3(_20235_),
    .A4(_09645_),
    .ZN(_09646_));
 NOR2_X1 _33420_ (.A1(_09614_),
    .A2(_09646_),
    .ZN(_20236_));
 INV_X1 _33421_ (.A(_20184_),
    .ZN(_09647_));
 INV_X1 _33422_ (.A(_20185_),
    .ZN(_09648_));
 BUF_X1 _33423_ (.A(_20187_),
    .Z(_09649_));
 INV_X1 _33424_ (.A(_20188_),
    .ZN(_09650_));
 INV_X1 _33425_ (.A(_20190_),
    .ZN(_09651_));
 INV_X1 _33426_ (.A(_20191_),
    .ZN(_09652_));
 BUF_X2 _33427_ (.A(_20195_),
    .Z(_09653_));
 AOI21_X2 _33428_ (.A(_20194_),
    .B1(_09653_),
    .B2(_20196_),
    .ZN(_09654_));
 INV_X1 _33429_ (.A(_09654_),
    .ZN(_09655_));
 BUF_X2 _33430_ (.A(_20193_),
    .Z(_09656_));
 AOI21_X1 _33431_ (.A(_20192_),
    .B1(_09655_),
    .B2(_09656_),
    .ZN(_09657_));
 OAI21_X1 _33432_ (.A(_09651_),
    .B1(_09652_),
    .B2(_09657_),
    .ZN(_09658_));
 BUF_X2 _33433_ (.A(_20199_),
    .Z(_09659_));
 AOI21_X2 _33434_ (.A(_20198_),
    .B1(_09659_),
    .B2(_20200_),
    .ZN(_09660_));
 NAND2_X1 _33435_ (.A1(_09659_),
    .A2(_09633_),
    .ZN(_09661_));
 OAI21_X1 _33436_ (.A(_09615_),
    .B1(_09641_),
    .B2(_09609_),
    .ZN(_09662_));
 AOI21_X1 _33437_ (.A(_20206_),
    .B1(_09594_),
    .B2(_09662_),
    .ZN(_09663_));
 OAI21_X1 _33438_ (.A(_09634_),
    .B1(_09663_),
    .B2(_09636_),
    .ZN(_09664_));
 AOI21_X1 _33439_ (.A(_20202_),
    .B1(_09590_),
    .B2(_09664_),
    .ZN(_09665_));
 OAI21_X1 _33440_ (.A(_09660_),
    .B1(_09661_),
    .B2(_09665_),
    .ZN(_09666_));
 INV_X1 _33441_ (.A(_09656_),
    .ZN(_09667_));
 BUF_X2 _33442_ (.A(_20197_),
    .Z(_09668_));
 NAND2_X2 _33443_ (.A1(_09653_),
    .A2(_09668_),
    .ZN(_09669_));
 NOR3_X2 _33444_ (.A1(_09652_),
    .A2(_09667_),
    .A3(_09669_),
    .ZN(_09670_));
 AOI21_X1 _33445_ (.A(_09658_),
    .B1(_09666_),
    .B2(_09670_),
    .ZN(_09671_));
 BUF_X2 _33446_ (.A(_20189_),
    .Z(_09672_));
 INV_X1 _33447_ (.A(_09672_),
    .ZN(_09673_));
 OAI21_X1 _33448_ (.A(_09650_),
    .B1(_09671_),
    .B2(_09673_),
    .ZN(_09674_));
 AOI21_X1 _33449_ (.A(_20186_),
    .B1(_09649_),
    .B2(_09674_),
    .ZN(_09675_));
 OAI21_X2 _33450_ (.A(_09647_),
    .B1(_09648_),
    .B2(_09675_),
    .ZN(_09676_));
 AOI21_X4 _33451_ (.A(_20182_),
    .B1(_20183_),
    .B2(_09676_),
    .ZN(_09677_));
 NOR4_X1 _33452_ (.A1(_09591_),
    .A2(_09609_),
    .A3(_09595_),
    .A4(_09661_),
    .ZN(_09678_));
 NOR2_X1 _33453_ (.A1(_09625_),
    .A2(_09642_),
    .ZN(_09679_));
 AOI21_X2 _33454_ (.A(_09666_),
    .B1(_09678_),
    .B2(_09679_),
    .ZN(_09680_));
 INV_X1 _33455_ (.A(_09680_),
    .ZN(_09681_));
 AOI21_X2 _33456_ (.A(_09658_),
    .B1(_09670_),
    .B2(_09681_),
    .ZN(_09682_));
 XNOR2_X2 _33457_ (.A(_09672_),
    .B(_09682_),
    .ZN(_09683_));
 INV_X1 _33458_ (.A(_20194_),
    .ZN(_09684_));
 AOI21_X1 _33459_ (.A(_20196_),
    .B1(_09668_),
    .B2(_20198_),
    .ZN(_09685_));
 NAND2_X1 _33460_ (.A1(_09668_),
    .A2(_09659_),
    .ZN(_09686_));
 AOI21_X1 _33461_ (.A(_20200_),
    .B1(_09633_),
    .B2(_20202_),
    .ZN(_09687_));
 OAI21_X1 _33462_ (.A(_09685_),
    .B1(_09686_),
    .B2(_09687_),
    .ZN(_09688_));
 NAND2_X1 _33463_ (.A1(_09633_),
    .A2(_09590_),
    .ZN(_09689_));
 INV_X1 _33464_ (.A(_20218_),
    .ZN(_09690_));
 OAI21_X1 _33465_ (.A(_09601_),
    .B1(_09690_),
    .B2(_09603_),
    .ZN(_09691_));
 AOI21_X1 _33466_ (.A(_09600_),
    .B1(_09691_),
    .B2(_09605_),
    .ZN(_09692_));
 OAI21_X1 _33467_ (.A(_09599_),
    .B1(_09692_),
    .B2(_09607_),
    .ZN(_09693_));
 AOI21_X1 _33468_ (.A(_09598_),
    .B1(_09612_),
    .B2(_09693_),
    .ZN(_09694_));
 NOR3_X1 _33469_ (.A1(_09686_),
    .A2(_09689_),
    .A3(_09694_),
    .ZN(_09695_));
 OAI21_X1 _33470_ (.A(_09653_),
    .B1(_09688_),
    .B2(_09695_),
    .ZN(_09696_));
 NAND2_X1 _33471_ (.A1(_09684_),
    .A2(_09696_),
    .ZN(_09697_));
 AOI21_X1 _33472_ (.A(_20192_),
    .B1(_09697_),
    .B2(_09656_),
    .ZN(_09698_));
 OAI21_X1 _33473_ (.A(_09651_),
    .B1(_09652_),
    .B2(_09698_),
    .ZN(_09699_));
 AOI21_X2 _33474_ (.A(_20188_),
    .B1(_09699_),
    .B2(_09672_),
    .ZN(_09700_));
 XNOR2_X2 _33475_ (.A(_09649_),
    .B(_09700_),
    .ZN(_09701_));
 OR2_X1 _33476_ (.A1(_09661_),
    .A2(_09669_),
    .ZN(_09702_));
 OAI221_X2 _33477_ (.A(_09654_),
    .B1(_09660_),
    .B2(_09669_),
    .C1(_09702_),
    .C2(_09644_),
    .ZN(_09703_));
 XNOR2_X2 _33478_ (.A(_09656_),
    .B(_09703_),
    .ZN(_09704_));
 XNOR2_X1 _33479_ (.A(_09590_),
    .B(_09613_),
    .ZN(_09705_));
 OAI21_X1 _33480_ (.A(_09687_),
    .B1(_09689_),
    .B2(_09593_),
    .ZN(_09706_));
 NOR2_X1 _33481_ (.A1(_09595_),
    .A2(_09689_),
    .ZN(_09707_));
 AOI21_X1 _33482_ (.A(_09706_),
    .B1(_09707_),
    .B2(_09617_),
    .ZN(_09708_));
 XNOR2_X1 _33483_ (.A(_09659_),
    .B(_09708_),
    .ZN(_09709_));
 NAND3_X1 _33484_ (.A1(_09705_),
    .A2(_20235_),
    .A3(_09709_),
    .ZN(_09710_));
 INV_X1 _33485_ (.A(_09653_),
    .ZN(_09711_));
 NOR3_X1 _33486_ (.A1(_09613_),
    .A2(_09686_),
    .A3(_09689_),
    .ZN(_09712_));
 NOR2_X1 _33487_ (.A1(_09688_),
    .A2(_09712_),
    .ZN(_09713_));
 XNOR2_X2 _33488_ (.A(_09711_),
    .B(_09713_),
    .ZN(_09714_));
 XOR2_X2 _33489_ (.A(_09668_),
    .B(_09680_),
    .Z(_09715_));
 OR3_X1 _33490_ (.A1(_09710_),
    .A2(_09714_),
    .A3(_09715_),
    .ZN(_09716_));
 OAI21_X1 _33491_ (.A(_09684_),
    .B1(_09711_),
    .B2(_09685_),
    .ZN(_09717_));
 AOI21_X1 _33492_ (.A(_20192_),
    .B1(_09717_),
    .B2(_09656_),
    .ZN(_09718_));
 NAND4_X1 _33493_ (.A1(_09656_),
    .A2(_09653_),
    .A3(_09668_),
    .A4(_09659_),
    .ZN(_09719_));
 OAI21_X1 _33494_ (.A(_09718_),
    .B1(_09719_),
    .B2(_09708_),
    .ZN(_09720_));
 XNOR2_X2 _33495_ (.A(_20191_),
    .B(_09720_),
    .ZN(_09721_));
 NOR3_X1 _33496_ (.A1(_09704_),
    .A2(_09716_),
    .A3(_09721_),
    .ZN(_09722_));
 NAND3_X1 _33497_ (.A1(_09683_),
    .A2(_09701_),
    .A3(_09722_),
    .ZN(_09723_));
 INV_X1 _33498_ (.A(_09600_),
    .ZN(_09724_));
 OAI21_X1 _33499_ (.A(_09599_),
    .B1(_09724_),
    .B2(_09607_),
    .ZN(_09725_));
 AOI21_X1 _33500_ (.A(_09596_),
    .B1(_09610_),
    .B2(_09725_),
    .ZN(_09726_));
 OAI21_X1 _33501_ (.A(_09615_),
    .B1(_09726_),
    .B2(_09609_),
    .ZN(_09727_));
 AOI21_X1 _33502_ (.A(_09706_),
    .B1(_09707_),
    .B2(_09727_),
    .ZN(_09728_));
 OAI21_X1 _33503_ (.A(_09718_),
    .B1(_09719_),
    .B2(_09728_),
    .ZN(_09729_));
 AOI21_X1 _33504_ (.A(_20190_),
    .B1(_20191_),
    .B2(_09729_),
    .ZN(_09730_));
 OAI21_X1 _33505_ (.A(_09650_),
    .B1(_09730_),
    .B2(_09673_),
    .ZN(_09731_));
 AOI21_X1 _33506_ (.A(_20186_),
    .B1(_09649_),
    .B2(_09731_),
    .ZN(_09732_));
 OAI21_X1 _33507_ (.A(_09647_),
    .B1(_09648_),
    .B2(_09732_),
    .ZN(_09733_));
 XNOR2_X2 _33508_ (.A(_20183_),
    .B(_09733_),
    .ZN(_09734_));
 INV_X1 _33509_ (.A(_20186_),
    .ZN(_09735_));
 INV_X1 _33510_ (.A(_09649_),
    .ZN(_09736_));
 AOI21_X1 _33511_ (.A(_09600_),
    .B1(_20216_),
    .B2(_09605_),
    .ZN(_09737_));
 OAI21_X1 _33512_ (.A(_09641_),
    .B1(_09642_),
    .B2(_09737_),
    .ZN(_09738_));
 AOI21_X1 _33513_ (.A(_09639_),
    .B1(_09640_),
    .B2(_09738_),
    .ZN(_09739_));
 OAI221_X1 _33514_ (.A(_09654_),
    .B1(_09660_),
    .B2(_09669_),
    .C1(_09702_),
    .C2(_09739_),
    .ZN(_09740_));
 AOI21_X1 _33515_ (.A(_20192_),
    .B1(_09740_),
    .B2(_09656_),
    .ZN(_09741_));
 OAI21_X1 _33516_ (.A(_09651_),
    .B1(_09652_),
    .B2(_09741_),
    .ZN(_09742_));
 AOI21_X1 _33517_ (.A(_20188_),
    .B1(_09742_),
    .B2(_09672_),
    .ZN(_09743_));
 OAI21_X1 _33518_ (.A(_09735_),
    .B1(_09736_),
    .B2(_09743_),
    .ZN(_09744_));
 XNOR2_X2 _33519_ (.A(_20185_),
    .B(_09744_),
    .ZN(_09745_));
 NOR3_X1 _33520_ (.A1(_09723_),
    .A2(_09734_),
    .A3(_09745_),
    .ZN(_09746_));
 XOR2_X1 _33521_ (.A(_09677_),
    .B(_09746_),
    .Z(_14450_));
 OR4_X1 _33522_ (.A1(\g_row[3].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09747_));
 OAI21_X2 _33523_ (.A(_07176_),
    .B1(_09747_),
    .B2(\g_row[3].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09748_));
 AND4_X1 _33524_ (.A1(\g_row[3].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09749_));
 AOI21_X4 _33525_ (.A(_07180_),
    .B1(_09749_),
    .B2(\g_row[3].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09750_));
 INV_X1 _33526_ (.A(_14448_),
    .ZN(_09751_));
 AOI21_X1 _33527_ (.A(_09748_),
    .B1(_09750_),
    .B2(_09751_),
    .ZN(_00401_));
 INV_X1 _33528_ (.A(_20225_),
    .ZN(_09752_));
 AOI21_X1 _33529_ (.A(_09748_),
    .B1(_09750_),
    .B2(_09752_),
    .ZN(_00402_));
 INV_X1 _33530_ (.A(_14456_),
    .ZN(_09753_));
 AOI21_X1 _33531_ (.A(_09748_),
    .B1(_09750_),
    .B2(_09753_),
    .ZN(_00403_));
 XOR2_X1 _33532_ (.A(_14455_),
    .B(_20234_),
    .Z(_09754_));
 AOI21_X1 _33533_ (.A(_09748_),
    .B1(_09750_),
    .B2(_09754_),
    .ZN(_00404_));
 AOI21_X1 _33534_ (.A(_20229_),
    .B1(_20230_),
    .B2(_20224_),
    .ZN(_09755_));
 INV_X1 _33535_ (.A(_09755_),
    .ZN(_09756_));
 AOI21_X1 _33536_ (.A(_20233_),
    .B1(_09756_),
    .B2(_20234_),
    .ZN(_09757_));
 XNOR2_X1 _33537_ (.A(\g_row[3].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20231_),
    .ZN(_09758_));
 XNOR2_X1 _33538_ (.A(_07174_),
    .B(_09758_),
    .ZN(_09759_));
 XNOR2_X1 _33539_ (.A(_09757_),
    .B(_09759_),
    .ZN(_09760_));
 AOI21_X1 _33540_ (.A(_09748_),
    .B1(_09750_),
    .B2(_09760_),
    .ZN(_00405_));
 INV_X1 _33541_ (.A(_09748_),
    .ZN(_09761_));
 NAND2_X4 _33542_ (.A1(_09761_),
    .A2(_09750_),
    .ZN(_09762_));
 INV_X1 _33543_ (.A(_14450_),
    .ZN(_14446_));
 NAND2_X1 _33544_ (.A1(_20238_),
    .A2(_14446_),
    .ZN(_09763_));
 NAND3_X1 _33545_ (.A1(_09705_),
    .A2(_09646_),
    .A3(_14450_),
    .ZN(_09764_));
 AOI21_X1 _33546_ (.A(_09762_),
    .B1(_09763_),
    .B2(_09764_),
    .ZN(_00400_));
 XNOR2_X1 _33547_ (.A(_20237_),
    .B(_09709_),
    .ZN(_09765_));
 INV_X1 _33548_ (.A(_20238_),
    .ZN(_09766_));
 MUX2_X1 _33549_ (.A(_09765_),
    .B(_09766_),
    .S(_14450_),
    .Z(_09767_));
 NOR2_X1 _33550_ (.A1(_09762_),
    .A2(_09767_),
    .ZN(_00406_));
 XNOR2_X1 _33551_ (.A(_09710_),
    .B(_09715_),
    .ZN(_09768_));
 MUX2_X1 _33552_ (.A(_09768_),
    .B(_09765_),
    .S(_14450_),
    .Z(_09769_));
 NOR2_X1 _33553_ (.A1(_09762_),
    .A2(_09769_),
    .ZN(_00407_));
 INV_X1 _33554_ (.A(_09715_),
    .ZN(_09770_));
 AND3_X1 _33555_ (.A1(_20237_),
    .A2(_09709_),
    .A3(_09770_),
    .ZN(_09771_));
 XOR2_X1 _33556_ (.A(_09714_),
    .B(_09771_),
    .Z(_09772_));
 MUX2_X1 _33557_ (.A(_09772_),
    .B(_09768_),
    .S(_14450_),
    .Z(_09773_));
 NOR2_X1 _33558_ (.A1(_09762_),
    .A2(_09773_),
    .ZN(_00408_));
 XNOR2_X1 _33559_ (.A(_09704_),
    .B(_09716_),
    .ZN(_09774_));
 MUX2_X1 _33560_ (.A(_09774_),
    .B(_09772_),
    .S(_14450_),
    .Z(_09775_));
 NOR2_X1 _33561_ (.A1(_09762_),
    .A2(_09775_),
    .ZN(_00409_));
 NOR2_X1 _33562_ (.A1(_09704_),
    .A2(_09714_),
    .ZN(_09776_));
 NAND2_X1 _33563_ (.A1(_09771_),
    .A2(_09776_),
    .ZN(_09777_));
 XNOR2_X1 _33564_ (.A(_09721_),
    .B(_09777_),
    .ZN(_09778_));
 MUX2_X1 _33565_ (.A(_09778_),
    .B(_09774_),
    .S(_14450_),
    .Z(_09779_));
 NOR2_X1 _33566_ (.A1(_09762_),
    .A2(_09779_),
    .ZN(_00410_));
 XNOR2_X1 _33567_ (.A(_09683_),
    .B(_09722_),
    .ZN(_09780_));
 MUX2_X1 _33568_ (.A(_09780_),
    .B(_09778_),
    .S(_14450_),
    .Z(_09781_));
 NOR2_X1 _33569_ (.A1(_09762_),
    .A2(_09781_),
    .ZN(_00411_));
 INV_X1 _33570_ (.A(_09683_),
    .ZN(_09782_));
 NOR3_X1 _33571_ (.A1(_09782_),
    .A2(_09721_),
    .A3(_09777_),
    .ZN(_09783_));
 XNOR2_X1 _33572_ (.A(_09701_),
    .B(_09783_),
    .ZN(_09784_));
 MUX2_X1 _33573_ (.A(_09784_),
    .B(_09780_),
    .S(_14450_),
    .Z(_09785_));
 NOR2_X1 _33574_ (.A1(_09762_),
    .A2(_09785_),
    .ZN(_00412_));
 NOR2_X1 _33575_ (.A1(_09723_),
    .A2(_09745_),
    .ZN(_09786_));
 AOI21_X1 _33576_ (.A(_09762_),
    .B1(_09784_),
    .B2(_09786_),
    .ZN(_09787_));
 AND2_X1 _33577_ (.A1(_09723_),
    .A2(_09745_),
    .ZN(_09788_));
 AOI21_X1 _33578_ (.A(_09788_),
    .B1(_09786_),
    .B2(_09734_),
    .ZN(_09789_));
 OAI21_X1 _33579_ (.A(_09787_),
    .B1(_09789_),
    .B2(_09677_),
    .ZN(_09790_));
 OR2_X1 _33580_ (.A1(_09746_),
    .A2(_09784_),
    .ZN(_09791_));
 AOI21_X1 _33581_ (.A(_09790_),
    .B1(_09791_),
    .B2(_09677_),
    .ZN(_00413_));
 INV_X1 _33582_ (.A(_09734_),
    .ZN(_09792_));
 NAND2_X1 _33583_ (.A1(_09701_),
    .A2(_09783_),
    .ZN(_09793_));
 AOI21_X1 _33584_ (.A(_09745_),
    .B1(_09793_),
    .B2(_09723_),
    .ZN(_09794_));
 NAND2_X1 _33585_ (.A1(_09792_),
    .A2(_09794_),
    .ZN(_09795_));
 OAI21_X1 _33586_ (.A(_09734_),
    .B1(_09745_),
    .B2(_09793_),
    .ZN(_09796_));
 NAND2_X1 _33587_ (.A1(_09795_),
    .A2(_09796_),
    .ZN(_09797_));
 AOI21_X1 _33588_ (.A(_09723_),
    .B1(_09792_),
    .B2(_09793_),
    .ZN(_09798_));
 MUX2_X1 _33589_ (.A(_09798_),
    .B(_09723_),
    .S(_09745_),
    .Z(_09799_));
 MUX2_X1 _33590_ (.A(_09797_),
    .B(_09799_),
    .S(_09677_),
    .Z(_09800_));
 NOR2_X1 _33591_ (.A1(_09762_),
    .A2(_09800_),
    .ZN(_00414_));
 CLKBUF_X2 _33592_ (.A(_20262_),
    .Z(_09801_));
 AOI21_X1 _33593_ (.A(_20261_),
    .B1(_09801_),
    .B2(_20263_),
    .ZN(_09802_));
 BUF_X1 _33594_ (.A(_20264_),
    .Z(_09803_));
 NAND2_X1 _33595_ (.A1(_09801_),
    .A2(_09803_),
    .ZN(_09804_));
 CLKBUF_X2 _33596_ (.A(_20267_),
    .Z(_09805_));
 AOI21_X1 _33597_ (.A(_20265_),
    .B1(_20266_),
    .B2(_09805_),
    .ZN(_09806_));
 OAI21_X1 _33598_ (.A(_09802_),
    .B1(_09804_),
    .B2(_09806_),
    .ZN(_09807_));
 INV_X1 _33599_ (.A(_20269_),
    .ZN(_09808_));
 CLKBUF_X2 _33600_ (.A(_20271_),
    .Z(_09809_));
 INV_X1 _33601_ (.A(_20273_),
    .ZN(_09810_));
 AOI21_X1 _33602_ (.A(_20275_),
    .B1(_20276_),
    .B2(_20277_),
    .ZN(_09811_));
 INV_X1 _33603_ (.A(_20274_),
    .ZN(_09812_));
 OAI21_X1 _33604_ (.A(_09810_),
    .B1(_09811_),
    .B2(_09812_),
    .ZN(_09813_));
 CLKBUF_X2 _33605_ (.A(_20272_),
    .Z(_09814_));
 AOI21_X1 _33606_ (.A(_09809_),
    .B1(_09813_),
    .B2(_09814_),
    .ZN(_09815_));
 INV_X1 _33607_ (.A(_20270_),
    .ZN(_09816_));
 OAI21_X1 _33608_ (.A(_09808_),
    .B1(_09815_),
    .B2(_09816_),
    .ZN(_09817_));
 INV_X1 _33609_ (.A(_20266_),
    .ZN(_09818_));
 CLKBUF_X2 _33610_ (.A(_20268_),
    .Z(_09819_));
 INV_X1 _33611_ (.A(_09819_),
    .ZN(_09820_));
 NOR3_X2 _33612_ (.A1(_09818_),
    .A2(_09820_),
    .A3(_09804_),
    .ZN(_09821_));
 AOI21_X2 _33613_ (.A(_09807_),
    .B1(_09817_),
    .B2(_09821_),
    .ZN(_09822_));
 XNOR2_X2 _33614_ (.A(_20260_),
    .B(_09822_),
    .ZN(_09823_));
 INV_X1 _33615_ (.A(_09823_),
    .ZN(_09824_));
 INV_X1 _33616_ (.A(_20265_),
    .ZN(_09825_));
 AOI21_X1 _33617_ (.A(_09805_),
    .B1(_09819_),
    .B2(_09817_),
    .ZN(_09826_));
 OAI21_X1 _33618_ (.A(_09825_),
    .B1(_09826_),
    .B2(_09818_),
    .ZN(_09827_));
 XNOR2_X1 _33619_ (.A(_09803_),
    .B(_09827_),
    .ZN(_09828_));
 XNOR2_X1 _33620_ (.A(_09820_),
    .B(_09817_),
    .ZN(_09829_));
 INV_X1 _33621_ (.A(_20259_),
    .ZN(_09830_));
 INV_X1 _33622_ (.A(_20260_),
    .ZN(_09831_));
 AOI21_X1 _33623_ (.A(_20263_),
    .B1(_09803_),
    .B2(_20265_),
    .ZN(_09832_));
 INV_X1 _33624_ (.A(_09832_),
    .ZN(_09833_));
 AOI21_X1 _33625_ (.A(_20261_),
    .B1(_09833_),
    .B2(_09801_),
    .ZN(_09834_));
 OAI21_X1 _33626_ (.A(_09830_),
    .B1(_09831_),
    .B2(_09834_),
    .ZN(_09835_));
 INV_X1 _33627_ (.A(_09801_),
    .ZN(_09836_));
 NAND2_X1 _33628_ (.A1(_09803_),
    .A2(_20266_),
    .ZN(_09837_));
 NOR3_X2 _33629_ (.A1(_09831_),
    .A2(_09836_),
    .A3(_09837_),
    .ZN(_09838_));
 AOI21_X2 _33630_ (.A(_09805_),
    .B1(_09819_),
    .B2(_20269_),
    .ZN(_09839_));
 OAI21_X1 _33631_ (.A(_09810_),
    .B1(_09812_),
    .B2(_14460_),
    .ZN(_09840_));
 AOI21_X2 _33632_ (.A(_09809_),
    .B1(_09840_),
    .B2(_09814_),
    .ZN(_09841_));
 NAND2_X1 _33633_ (.A1(_09819_),
    .A2(_20270_),
    .ZN(_09842_));
 NOR2_X1 _33634_ (.A1(_09841_),
    .A2(_09842_),
    .ZN(_09843_));
 INV_X1 _33635_ (.A(_09843_),
    .ZN(_09844_));
 NAND2_X1 _33636_ (.A1(_09839_),
    .A2(_09844_),
    .ZN(_09845_));
 AOI21_X2 _33637_ (.A(_09835_),
    .B1(_09838_),
    .B2(_09845_),
    .ZN(_09846_));
 XNOR2_X2 _33638_ (.A(_20258_),
    .B(_09846_),
    .ZN(_20292_));
 AOI21_X1 _33639_ (.A(_09820_),
    .B1(_09816_),
    .B2(_09808_),
    .ZN(_09847_));
 NOR2_X1 _33640_ (.A1(_09805_),
    .A2(_09847_),
    .ZN(_09848_));
 XNOR2_X1 _33641_ (.A(_09818_),
    .B(_09848_),
    .ZN(_09849_));
 XNOR2_X1 _33642_ (.A(_14460_),
    .B(_20274_),
    .ZN(_09850_));
 NOR4_X1 _33643_ (.A1(_14461_),
    .A2(\g_row[3].g_col[2].mult.adder.a[0] ),
    .A3(_20278_),
    .A4(_09850_),
    .ZN(_09851_));
 XNOR2_X1 _33644_ (.A(_09816_),
    .B(_09841_),
    .ZN(_09852_));
 XNOR2_X1 _33645_ (.A(_09814_),
    .B(_09813_),
    .ZN(_09853_));
 NAND4_X1 _33646_ (.A1(_09849_),
    .A2(_09851_),
    .A3(_09852_),
    .A4(_09853_),
    .ZN(_09854_));
 OAI21_X1 _33647_ (.A(_09832_),
    .B1(_09837_),
    .B2(_09839_),
    .ZN(_09855_));
 NOR2_X1 _33648_ (.A1(_09837_),
    .A2(_09844_),
    .ZN(_09856_));
 NOR2_X1 _33649_ (.A1(_09855_),
    .A2(_09856_),
    .ZN(_09857_));
 XNOR2_X1 _33650_ (.A(_09801_),
    .B(_09857_),
    .ZN(_09858_));
 NOR4_X1 _33651_ (.A1(_09829_),
    .A2(_20292_),
    .A3(_09854_),
    .A4(_09858_),
    .ZN(_09859_));
 AND2_X1 _33652_ (.A1(_09828_),
    .A2(_09859_),
    .ZN(_09860_));
 NOR2_X1 _33653_ (.A1(_09824_),
    .A2(_09860_),
    .ZN(_20293_));
 INV_X1 _33654_ (.A(_20239_),
    .ZN(_09861_));
 INV_X1 _33655_ (.A(_20240_),
    .ZN(_09862_));
 INV_X1 _33656_ (.A(_20243_),
    .ZN(_09863_));
 INV_X1 _33657_ (.A(_20244_),
    .ZN(_09864_));
 INV_X1 _33658_ (.A(_20249_),
    .ZN(_09865_));
 CLKBUF_X3 _33659_ (.A(_20252_),
    .Z(_09866_));
 AOI21_X2 _33660_ (.A(_20251_),
    .B1(_09866_),
    .B2(_20253_),
    .ZN(_09867_));
 CLKBUF_X2 _33661_ (.A(_20250_),
    .Z(_09868_));
 INV_X1 _33662_ (.A(_09868_),
    .ZN(_09869_));
 OAI21_X1 _33663_ (.A(_09865_),
    .B1(_09867_),
    .B2(_09869_),
    .ZN(_09870_));
 AOI21_X1 _33664_ (.A(_20247_),
    .B1(_20248_),
    .B2(_09870_),
    .ZN(_09871_));
 BUF_X2 _33665_ (.A(_20256_),
    .Z(_09872_));
 AND2_X1 _33666_ (.A1(_09872_),
    .A2(_20258_),
    .ZN(_09873_));
 AOI21_X1 _33667_ (.A(_20261_),
    .B1(_09855_),
    .B2(_09801_),
    .ZN(_09874_));
 OAI21_X1 _33668_ (.A(_09830_),
    .B1(_09831_),
    .B2(_09874_),
    .ZN(_09875_));
 AOI221_X2 _33669_ (.A(_20255_),
    .B1(_09872_),
    .B2(_20257_),
    .C1(_09873_),
    .C2(_09875_),
    .ZN(_09876_));
 BUF_X2 _33670_ (.A(_20254_),
    .Z(_09877_));
 NAND4_X1 _33671_ (.A1(_20248_),
    .A2(_09868_),
    .A3(_09866_),
    .A4(_09877_),
    .ZN(_09878_));
 OAI21_X1 _33672_ (.A(_09871_),
    .B1(_09876_),
    .B2(_09878_),
    .ZN(_09879_));
 BUF_X2 _33673_ (.A(_20246_),
    .Z(_09880_));
 AOI21_X1 _33674_ (.A(_20245_),
    .B1(_09879_),
    .B2(_09880_),
    .ZN(_09881_));
 OAI21_X1 _33675_ (.A(_09863_),
    .B1(_09864_),
    .B2(_09881_),
    .ZN(_09882_));
 AOI21_X2 _33676_ (.A(_20241_),
    .B1(_20242_),
    .B2(_09882_),
    .ZN(_09883_));
 OAI21_X4 _33677_ (.A(_09861_),
    .B1(_09862_),
    .B2(_09883_),
    .ZN(_09884_));
 INV_X1 _33678_ (.A(_20251_),
    .ZN(_09885_));
 INV_X1 _33679_ (.A(_09866_),
    .ZN(_09886_));
 AOI21_X1 _33680_ (.A(_20253_),
    .B1(_09877_),
    .B2(_20255_),
    .ZN(_09887_));
 OAI21_X1 _33681_ (.A(_09885_),
    .B1(_09886_),
    .B2(_09887_),
    .ZN(_09888_));
 AOI21_X1 _33682_ (.A(_20249_),
    .B1(_09888_),
    .B2(_09868_),
    .ZN(_09889_));
 NAND4_X1 _33683_ (.A1(_09868_),
    .A2(_09866_),
    .A3(_09877_),
    .A4(_09872_),
    .ZN(_09890_));
 AOI21_X1 _33684_ (.A(_20257_),
    .B1(_20258_),
    .B2(_20259_),
    .ZN(_09891_));
 NAND2_X1 _33685_ (.A1(_20258_),
    .A2(_20260_),
    .ZN(_09892_));
 OAI21_X1 _33686_ (.A(_09891_),
    .B1(_09892_),
    .B2(_09802_),
    .ZN(_09893_));
 NOR2_X1 _33687_ (.A1(_09804_),
    .A2(_09892_),
    .ZN(_09894_));
 INV_X1 _33688_ (.A(_09809_),
    .ZN(_09895_));
 OAI21_X1 _33689_ (.A(_09808_),
    .B1(_09895_),
    .B2(_09816_),
    .ZN(_09896_));
 AOI21_X1 _33690_ (.A(_09805_),
    .B1(_09819_),
    .B2(_09896_),
    .ZN(_09897_));
 OAI21_X1 _33691_ (.A(_09825_),
    .B1(_09897_),
    .B2(_09818_),
    .ZN(_09898_));
 AOI21_X1 _33692_ (.A(_09893_),
    .B1(_09894_),
    .B2(_09898_),
    .ZN(_09899_));
 OAI21_X1 _33693_ (.A(_09889_),
    .B1(_09890_),
    .B2(_09899_),
    .ZN(_09900_));
 AOI21_X1 _33694_ (.A(_20247_),
    .B1(_20248_),
    .B2(_09900_),
    .ZN(_09901_));
 INV_X1 _33695_ (.A(_09901_),
    .ZN(_09902_));
 AOI21_X1 _33696_ (.A(_20245_),
    .B1(_09902_),
    .B2(_09880_),
    .ZN(_09903_));
 OAI21_X1 _33697_ (.A(_09863_),
    .B1(_09864_),
    .B2(_09903_),
    .ZN(_09904_));
 AOI21_X2 _33698_ (.A(_20241_),
    .B1(_20242_),
    .B2(_09904_),
    .ZN(_09905_));
 XNOR2_X2 _33699_ (.A(_20240_),
    .B(_09905_),
    .ZN(_09906_));
 INV_X1 _33700_ (.A(_09906_),
    .ZN(_09907_));
 INV_X1 _33701_ (.A(_20247_),
    .ZN(_09908_));
 INV_X1 _33702_ (.A(_20248_),
    .ZN(_09909_));
 AOI21_X2 _33703_ (.A(_20255_),
    .B1(_09872_),
    .B2(_20257_),
    .ZN(_09910_));
 NAND2_X1 _33704_ (.A1(_09866_),
    .A2(_09877_),
    .ZN(_09911_));
 NAND3_X1 _33705_ (.A1(_09866_),
    .A2(_09877_),
    .A3(_09873_),
    .ZN(_09912_));
 AOI21_X1 _33706_ (.A(_09809_),
    .B1(_20273_),
    .B2(_09814_),
    .ZN(_09913_));
 OAI21_X1 _33707_ (.A(_09839_),
    .B1(_09842_),
    .B2(_09913_),
    .ZN(_09914_));
 AOI21_X1 _33708_ (.A(_09835_),
    .B1(_09838_),
    .B2(_09914_),
    .ZN(_09915_));
 OAI221_X1 _33709_ (.A(_09867_),
    .B1(_09910_),
    .B2(_09911_),
    .C1(_09912_),
    .C2(_09915_),
    .ZN(_09916_));
 AOI21_X1 _33710_ (.A(_20249_),
    .B1(_09916_),
    .B2(_09868_),
    .ZN(_09917_));
 OAI21_X1 _33711_ (.A(_09908_),
    .B1(_09909_),
    .B2(_09917_),
    .ZN(_09918_));
 AOI21_X1 _33712_ (.A(_20245_),
    .B1(_09918_),
    .B2(_09880_),
    .ZN(_09919_));
 OAI21_X1 _33713_ (.A(_09863_),
    .B1(_09864_),
    .B2(_09919_),
    .ZN(_09920_));
 XNOR2_X2 _33714_ (.A(_20242_),
    .B(_09920_),
    .ZN(_09921_));
 NAND2_X1 _33715_ (.A1(_09838_),
    .A2(_09873_),
    .ZN(_09922_));
 OAI21_X2 _33716_ (.A(_09876_),
    .B1(_09922_),
    .B2(_09844_),
    .ZN(_09923_));
 INV_X1 _33717_ (.A(_09923_),
    .ZN(_09924_));
 OAI21_X1 _33718_ (.A(_09871_),
    .B1(_09878_),
    .B2(_09924_),
    .ZN(_09925_));
 XOR2_X2 _33719_ (.A(_09880_),
    .B(_09925_),
    .Z(_09926_));
 NAND2_X1 _33720_ (.A1(_09877_),
    .A2(_09872_),
    .ZN(_09927_));
 OAI21_X1 _33721_ (.A(_09887_),
    .B1(_09927_),
    .B2(_09891_),
    .ZN(_09928_));
 INV_X1 _33722_ (.A(_20275_),
    .ZN(_09929_));
 OAI21_X1 _33723_ (.A(_09810_),
    .B1(_09929_),
    .B2(_09812_),
    .ZN(_09930_));
 AOI21_X1 _33724_ (.A(_09809_),
    .B1(_09930_),
    .B2(_09814_),
    .ZN(_09931_));
 OAI21_X1 _33725_ (.A(_09808_),
    .B1(_09931_),
    .B2(_09816_),
    .ZN(_09932_));
 AOI21_X1 _33726_ (.A(_09807_),
    .B1(_09821_),
    .B2(_09932_),
    .ZN(_09933_));
 NOR3_X1 _33727_ (.A1(_09927_),
    .A2(_09892_),
    .A3(_09933_),
    .ZN(_09934_));
 OAI21_X1 _33728_ (.A(_09866_),
    .B1(_09928_),
    .B2(_09934_),
    .ZN(_09935_));
 NAND2_X1 _33729_ (.A1(_09885_),
    .A2(_09935_),
    .ZN(_09936_));
 AOI21_X1 _33730_ (.A(_20249_),
    .B1(_09936_),
    .B2(_09868_),
    .ZN(_09937_));
 OAI21_X1 _33731_ (.A(_09908_),
    .B1(_09909_),
    .B2(_09937_),
    .ZN(_09938_));
 AOI21_X2 _33732_ (.A(_20245_),
    .B1(_09938_),
    .B2(_09880_),
    .ZN(_09939_));
 XNOR2_X2 _33733_ (.A(_20244_),
    .B(_09939_),
    .ZN(_09940_));
 OAI221_X2 _33734_ (.A(_09867_),
    .B1(_09910_),
    .B2(_09911_),
    .C1(_09912_),
    .C2(_09846_),
    .ZN(_09941_));
 XNOR2_X2 _33735_ (.A(_09869_),
    .B(_09941_),
    .ZN(_09942_));
 AOI21_X1 _33736_ (.A(_09893_),
    .B1(_09894_),
    .B2(_09827_),
    .ZN(_09943_));
 XNOR2_X1 _33737_ (.A(_09872_),
    .B(_09943_),
    .ZN(_09944_));
 AND3_X1 _33738_ (.A1(_09823_),
    .A2(_20292_),
    .A3(_09944_),
    .ZN(_09945_));
 NOR3_X1 _33739_ (.A1(_09822_),
    .A2(_09927_),
    .A3(_09892_),
    .ZN(_09946_));
 NOR2_X1 _33740_ (.A1(_09928_),
    .A2(_09946_),
    .ZN(_09947_));
 XNOR2_X2 _33741_ (.A(_09866_),
    .B(_09947_),
    .ZN(_09948_));
 XOR2_X2 _33742_ (.A(_09877_),
    .B(_09923_),
    .Z(_09949_));
 AND3_X1 _33743_ (.A1(_09945_),
    .A2(_09948_),
    .A3(_09949_),
    .ZN(_09950_));
 OAI21_X1 _33744_ (.A(_09889_),
    .B1(_09890_),
    .B2(_09943_),
    .ZN(_09951_));
 XNOR2_X2 _33745_ (.A(_09909_),
    .B(_09951_),
    .ZN(_09952_));
 AND3_X1 _33746_ (.A1(_09942_),
    .A2(_09950_),
    .A3(_09952_),
    .ZN(_09953_));
 NAND3_X1 _33747_ (.A1(_09926_),
    .A2(_09940_),
    .A3(_09953_),
    .ZN(_09954_));
 OR3_X1 _33748_ (.A1(_09907_),
    .A2(_09921_),
    .A3(_09954_),
    .ZN(_09955_));
 XNOR2_X1 _33749_ (.A(_09884_),
    .B(_09955_),
    .ZN(_09956_));
 BUF_X1 _33750_ (.A(_09956_),
    .Z(_14463_));
 INV_X1 _33751_ (.A(_14463_),
    .ZN(_14466_));
 OR4_X2 _33752_ (.A1(\g_row[3].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09957_));
 OAI21_X4 _33753_ (.A(_07394_),
    .B1(_09957_),
    .B2(\g_row[3].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09958_));
 AND4_X1 _33754_ (.A1(\g_row[3].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_09959_));
 AOI21_X4 _33755_ (.A(_07398_),
    .B1(_09959_),
    .B2(\g_row[3].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_09960_));
 INV_X1 _33756_ (.A(_14465_),
    .ZN(_09961_));
 AOI21_X1 _33757_ (.A(_09958_),
    .B1(_09960_),
    .B2(_09961_),
    .ZN(_00417_));
 INV_X1 _33758_ (.A(_20282_),
    .ZN(_09962_));
 AOI21_X1 _33759_ (.A(_09958_),
    .B1(_09960_),
    .B2(_09962_),
    .ZN(_00418_));
 INV_X1 _33760_ (.A(_14473_),
    .ZN(_09963_));
 AOI21_X1 _33761_ (.A(_09958_),
    .B1(_09960_),
    .B2(_09963_),
    .ZN(_00419_));
 XOR2_X2 _33762_ (.A(_14472_),
    .B(_20291_),
    .Z(_09964_));
 AOI21_X1 _33763_ (.A(_09958_),
    .B1(_09960_),
    .B2(_09964_),
    .ZN(_00420_));
 AOI21_X1 _33764_ (.A(_20286_),
    .B1(_20287_),
    .B2(_20281_),
    .ZN(_09965_));
 INV_X1 _33765_ (.A(_09965_),
    .ZN(_09966_));
 AOI21_X1 _33766_ (.A(_20290_),
    .B1(_09966_),
    .B2(_20291_),
    .ZN(_09967_));
 XNOR2_X1 _33767_ (.A(\g_row[3].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20288_),
    .ZN(_09968_));
 XNOR2_X1 _33768_ (.A(_07392_),
    .B(_09968_),
    .ZN(_09969_));
 XNOR2_X1 _33769_ (.A(_09967_),
    .B(_09969_),
    .ZN(_09970_));
 AOI21_X1 _33770_ (.A(_09958_),
    .B1(_09960_),
    .B2(_09970_),
    .ZN(_00421_));
 INV_X1 _33771_ (.A(_09958_),
    .ZN(_09971_));
 NAND2_X4 _33772_ (.A1(_09971_),
    .A2(_09960_),
    .ZN(_09972_));
 NAND2_X1 _33773_ (.A1(_20295_),
    .A2(_14463_),
    .ZN(_09973_));
 NAND3_X1 _33774_ (.A1(_09823_),
    .A2(_09860_),
    .A3(_14466_),
    .ZN(_09974_));
 AOI21_X2 _33775_ (.A(_09972_),
    .B1(_09973_),
    .B2(_09974_),
    .ZN(_00416_));
 INV_X1 _33776_ (.A(_20295_),
    .ZN(_09975_));
 XNOR2_X2 _33777_ (.A(_20294_),
    .B(_09944_),
    .ZN(_09976_));
 MUX2_X1 _33778_ (.A(_09975_),
    .B(_09976_),
    .S(_14463_),
    .Z(_09977_));
 NOR2_X1 _33779_ (.A1(_09972_),
    .A2(_09977_),
    .ZN(_00422_));
 XNOR2_X2 _33780_ (.A(_09945_),
    .B(_09949_),
    .ZN(_09978_));
 MUX2_X1 _33781_ (.A(_09976_),
    .B(_09978_),
    .S(_14463_),
    .Z(_09979_));
 NOR2_X1 _33782_ (.A1(_09972_),
    .A2(_09979_),
    .ZN(_00423_));
 AND3_X1 _33783_ (.A1(_20294_),
    .A2(_09944_),
    .A3(_09949_),
    .ZN(_09980_));
 XNOR2_X2 _33784_ (.A(_09948_),
    .B(_09980_),
    .ZN(_09981_));
 MUX2_X1 _33785_ (.A(_09978_),
    .B(_09981_),
    .S(_14463_),
    .Z(_09982_));
 NOR2_X1 _33786_ (.A1(_09972_),
    .A2(_09982_),
    .ZN(_00424_));
 XNOR2_X2 _33787_ (.A(_09942_),
    .B(_09950_),
    .ZN(_09983_));
 MUX2_X1 _33788_ (.A(_09981_),
    .B(_09983_),
    .S(_14463_),
    .Z(_09984_));
 NOR2_X1 _33789_ (.A1(_09972_),
    .A2(_09984_),
    .ZN(_00425_));
 AND3_X1 _33790_ (.A1(_09942_),
    .A2(_09948_),
    .A3(_09980_),
    .ZN(_09985_));
 XNOR2_X2 _33791_ (.A(_09952_),
    .B(_09985_),
    .ZN(_09986_));
 MUX2_X1 _33792_ (.A(_09983_),
    .B(_09986_),
    .S(_14463_),
    .Z(_09987_));
 NOR2_X1 _33793_ (.A1(_09972_),
    .A2(_09987_),
    .ZN(_00426_));
 XNOR2_X2 _33794_ (.A(_09926_),
    .B(_09953_),
    .ZN(_09988_));
 MUX2_X1 _33795_ (.A(_09986_),
    .B(_09988_),
    .S(_09956_),
    .Z(_09989_));
 NOR2_X1 _33796_ (.A1(_09972_),
    .A2(_09989_),
    .ZN(_00427_));
 NAND3_X2 _33797_ (.A1(_09926_),
    .A2(_09952_),
    .A3(_09985_),
    .ZN(_09990_));
 XNOR2_X1 _33798_ (.A(_09940_),
    .B(_09990_),
    .ZN(_09991_));
 NAND2_X1 _33799_ (.A1(_14463_),
    .A2(_09991_),
    .ZN(_09992_));
 OR2_X1 _33800_ (.A1(_14463_),
    .A2(_09988_),
    .ZN(_09993_));
 AOI21_X2 _33801_ (.A(_09972_),
    .B1(_09992_),
    .B2(_09993_),
    .ZN(_00428_));
 AND4_X1 _33802_ (.A1(_09940_),
    .A2(_09942_),
    .A3(_09950_),
    .A4(_09952_),
    .ZN(_09994_));
 AND2_X1 _33803_ (.A1(_09926_),
    .A2(_09994_),
    .ZN(_09995_));
 XNOR2_X2 _33804_ (.A(_09995_),
    .B(_09921_),
    .ZN(_09996_));
 NAND2_X1 _33805_ (.A1(_09921_),
    .A2(_09954_),
    .ZN(_09997_));
 NAND3_X1 _33806_ (.A1(_09884_),
    .A2(_09906_),
    .A3(_09997_),
    .ZN(_09998_));
 INV_X1 _33807_ (.A(_09955_),
    .ZN(_09999_));
 OAI21_X2 _33808_ (.A(_09998_),
    .B1(_09999_),
    .B2(_09884_),
    .ZN(_10000_));
 AOI22_X4 _33809_ (.A1(_09884_),
    .A2(_09996_),
    .B1(_10000_),
    .B2(_09991_),
    .ZN(_10001_));
 NOR2_X1 _33810_ (.A1(_09972_),
    .A2(_10001_),
    .ZN(_00429_));
 INV_X1 _33811_ (.A(_09940_),
    .ZN(_10002_));
 NOR2_X1 _33812_ (.A1(_10002_),
    .A2(_09990_),
    .ZN(_10003_));
 OAI21_X1 _33813_ (.A(_09995_),
    .B1(_09907_),
    .B2(_10003_),
    .ZN(_10004_));
 OAI21_X1 _33814_ (.A(_09997_),
    .B1(_10004_),
    .B2(_09921_),
    .ZN(_10005_));
 NOR2_X1 _33815_ (.A1(_09884_),
    .A2(_10005_),
    .ZN(_10006_));
 INV_X1 _33816_ (.A(_09921_),
    .ZN(_10007_));
 OAI21_X1 _33817_ (.A(_10007_),
    .B1(_10003_),
    .B2(_09995_),
    .ZN(_10008_));
 NOR2_X1 _33818_ (.A1(_09907_),
    .A2(_10008_),
    .ZN(_10009_));
 AOI21_X1 _33819_ (.A(_09906_),
    .B1(_10007_),
    .B2(_10003_),
    .ZN(_10010_));
 NOR2_X1 _33820_ (.A1(_10009_),
    .A2(_10010_),
    .ZN(_10011_));
 AOI21_X1 _33821_ (.A(_10006_),
    .B1(_10011_),
    .B2(_09884_),
    .ZN(_10012_));
 NOR2_X1 _33822_ (.A1(_09972_),
    .A2(_10012_),
    .ZN(_00430_));
 BUF_X2 _33823_ (.A(_20319_),
    .Z(_10013_));
 AOI21_X2 _33824_ (.A(_20318_),
    .B1(_10013_),
    .B2(_20320_),
    .ZN(_10014_));
 BUF_X2 _33825_ (.A(_20321_),
    .Z(_10015_));
 NAND2_X1 _33826_ (.A1(_10013_),
    .A2(_10015_),
    .ZN(_10016_));
 CLKBUF_X2 _33827_ (.A(_20324_),
    .Z(_10017_));
 AOI21_X1 _33828_ (.A(_20322_),
    .B1(_20323_),
    .B2(_10017_),
    .ZN(_10018_));
 OAI21_X1 _33829_ (.A(_10014_),
    .B1(_10016_),
    .B2(_10018_),
    .ZN(_10019_));
 INV_X1 _33830_ (.A(_20326_),
    .ZN(_10020_));
 CLKBUF_X2 _33831_ (.A(_20328_),
    .Z(_10021_));
 INV_X1 _33832_ (.A(_20330_),
    .ZN(_10022_));
 AOI21_X1 _33833_ (.A(_20332_),
    .B1(_20333_),
    .B2(_20334_),
    .ZN(_10023_));
 INV_X1 _33834_ (.A(_20331_),
    .ZN(_10024_));
 OAI21_X1 _33835_ (.A(_10022_),
    .B1(_10023_),
    .B2(_10024_),
    .ZN(_10025_));
 AOI21_X1 _33836_ (.A(_10021_),
    .B1(_10025_),
    .B2(_20329_),
    .ZN(_10026_));
 CLKBUF_X2 _33837_ (.A(_20327_),
    .Z(_10027_));
 INV_X1 _33838_ (.A(_10027_),
    .ZN(_10028_));
 OAI21_X2 _33839_ (.A(_10020_),
    .B1(_10026_),
    .B2(_10028_),
    .ZN(_10029_));
 INV_X1 _33840_ (.A(_20323_),
    .ZN(_10030_));
 BUF_X2 _33841_ (.A(_20325_),
    .Z(_10031_));
 INV_X1 _33842_ (.A(_10031_),
    .ZN(_10032_));
 NOR3_X1 _33843_ (.A1(_10030_),
    .A2(_10032_),
    .A3(_10016_),
    .ZN(_10033_));
 AOI21_X2 _33844_ (.A(_10019_),
    .B1(_10029_),
    .B2(_10033_),
    .ZN(_10034_));
 XNOR2_X2 _33845_ (.A(_20317_),
    .B(_10034_),
    .ZN(_10035_));
 INV_X1 _33846_ (.A(_10035_),
    .ZN(_10036_));
 INV_X1 _33847_ (.A(_20322_),
    .ZN(_10037_));
 AOI21_X1 _33848_ (.A(_10017_),
    .B1(_10031_),
    .B2(_10029_),
    .ZN(_10038_));
 OAI21_X2 _33849_ (.A(_10037_),
    .B1(_10038_),
    .B2(_10030_),
    .ZN(_10039_));
 XOR2_X2 _33850_ (.A(_10015_),
    .B(_10039_),
    .Z(_10040_));
 XNOR2_X2 _33851_ (.A(_10032_),
    .B(_10029_),
    .ZN(_10041_));
 CLKBUF_X3 _33852_ (.A(_20315_),
    .Z(_10042_));
 INV_X1 _33853_ (.A(_20316_),
    .ZN(_10043_));
 INV_X1 _33854_ (.A(_20317_),
    .ZN(_10044_));
 AOI21_X1 _33855_ (.A(_20320_),
    .B1(_10015_),
    .B2(_20322_),
    .ZN(_10045_));
 INV_X1 _33856_ (.A(_10045_),
    .ZN(_10046_));
 AOI21_X1 _33857_ (.A(_20318_),
    .B1(_10046_),
    .B2(_10013_),
    .ZN(_10047_));
 OAI21_X1 _33858_ (.A(_10043_),
    .B1(_10044_),
    .B2(_10047_),
    .ZN(_10048_));
 INV_X1 _33859_ (.A(_10013_),
    .ZN(_10049_));
 NAND2_X1 _33860_ (.A1(_10015_),
    .A2(_20323_),
    .ZN(_10050_));
 NOR3_X2 _33861_ (.A1(_10044_),
    .A2(_10049_),
    .A3(_10050_),
    .ZN(_10051_));
 AOI21_X2 _33862_ (.A(_10017_),
    .B1(_10031_),
    .B2(_20326_),
    .ZN(_10052_));
 OAI21_X1 _33863_ (.A(_10022_),
    .B1(_10024_),
    .B2(_14477_),
    .ZN(_10053_));
 AOI21_X1 _33864_ (.A(_10021_),
    .B1(_10053_),
    .B2(_20329_),
    .ZN(_10054_));
 NAND2_X1 _33865_ (.A1(_10031_),
    .A2(_10027_),
    .ZN(_10055_));
 NOR2_X1 _33866_ (.A1(_10054_),
    .A2(_10055_),
    .ZN(_10056_));
 INV_X1 _33867_ (.A(_10056_),
    .ZN(_10057_));
 NAND2_X1 _33868_ (.A1(_10052_),
    .A2(_10057_),
    .ZN(_10058_));
 AOI21_X1 _33869_ (.A(_10048_),
    .B1(_10051_),
    .B2(_10058_),
    .ZN(_10059_));
 XNOR2_X1 _33870_ (.A(_10042_),
    .B(_10059_),
    .ZN(_20349_));
 XNOR2_X1 _33871_ (.A(_10027_),
    .B(_10054_),
    .ZN(_10060_));
 INV_X1 _33872_ (.A(_20329_),
    .ZN(_10061_));
 XNOR2_X1 _33873_ (.A(_10061_),
    .B(_10025_),
    .ZN(_10062_));
 NOR2_X1 _33874_ (.A1(_10060_),
    .A2(_10062_),
    .ZN(_10063_));
 AOI21_X1 _33875_ (.A(_10032_),
    .B1(_10028_),
    .B2(_10020_),
    .ZN(_10064_));
 NOR2_X1 _33876_ (.A1(_10017_),
    .A2(_10064_),
    .ZN(_10065_));
 XNOR2_X1 _33877_ (.A(_10030_),
    .B(_10065_),
    .ZN(_10066_));
 XNOR2_X1 _33878_ (.A(_14477_),
    .B(_20331_),
    .ZN(_10067_));
 NOR4_X2 _33879_ (.A1(_14478_),
    .A2(\g_row[3].g_col[3].mult.adder.a[0] ),
    .A3(_20335_),
    .A4(_10067_),
    .ZN(_10068_));
 OAI21_X1 _33880_ (.A(_10045_),
    .B1(_10050_),
    .B2(_10052_),
    .ZN(_10069_));
 NOR2_X1 _33881_ (.A1(_10050_),
    .A2(_10057_),
    .ZN(_10070_));
 NOR2_X1 _33882_ (.A1(_10069_),
    .A2(_10070_),
    .ZN(_10071_));
 XNOR2_X1 _33883_ (.A(_10049_),
    .B(_10071_),
    .ZN(_10072_));
 NAND4_X2 _33884_ (.A1(_10063_),
    .A2(_10066_),
    .A3(_10068_),
    .A4(_10072_),
    .ZN(_10073_));
 NOR4_X4 _33885_ (.A1(_10040_),
    .A2(_10041_),
    .A3(_20349_),
    .A4(_10073_),
    .ZN(_10074_));
 NOR2_X1 _33886_ (.A1(_10036_),
    .A2(_10074_),
    .ZN(_20350_));
 INV_X1 _33887_ (.A(_20298_),
    .ZN(_10075_));
 INV_X1 _33888_ (.A(_20299_),
    .ZN(_10076_));
 CLKBUF_X2 _33889_ (.A(_20301_),
    .Z(_10077_));
 INV_X1 _33890_ (.A(_20302_),
    .ZN(_10078_));
 INV_X1 _33891_ (.A(_20304_),
    .ZN(_10079_));
 BUF_X1 _33892_ (.A(_20305_),
    .Z(_10080_));
 INV_X1 _33893_ (.A(_10080_),
    .ZN(_10081_));
 BUF_X2 _33894_ (.A(_20309_),
    .Z(_10082_));
 AOI21_X2 _33895_ (.A(_20308_),
    .B1(_10082_),
    .B2(_20310_),
    .ZN(_10083_));
 INV_X1 _33896_ (.A(_10083_),
    .ZN(_10084_));
 CLKBUF_X2 _33897_ (.A(_20307_),
    .Z(_10085_));
 AOI21_X1 _33898_ (.A(_20306_),
    .B1(_10084_),
    .B2(_10085_),
    .ZN(_10086_));
 OAI21_X1 _33899_ (.A(_10079_),
    .B1(_10081_),
    .B2(_10086_),
    .ZN(_10087_));
 INV_X1 _33900_ (.A(_10085_),
    .ZN(_10088_));
 BUF_X2 _33901_ (.A(_20311_),
    .Z(_10089_));
 NAND2_X2 _33902_ (.A1(_10082_),
    .A2(_10089_),
    .ZN(_10090_));
 NOR3_X2 _33903_ (.A1(_10081_),
    .A2(_10088_),
    .A3(_10090_),
    .ZN(_10091_));
 INV_X1 _33904_ (.A(_20312_),
    .ZN(_10092_));
 CLKBUF_X3 _33905_ (.A(_20313_),
    .Z(_10093_));
 INV_X1 _33906_ (.A(_10093_),
    .ZN(_10094_));
 BUF_X2 _33907_ (.A(_20314_),
    .Z(_10095_));
 AOI21_X1 _33908_ (.A(_20318_),
    .B1(_10069_),
    .B2(_10013_),
    .ZN(_10096_));
 OAI21_X1 _33909_ (.A(_10043_),
    .B1(_10044_),
    .B2(_10096_),
    .ZN(_10097_));
 AOI21_X1 _33910_ (.A(_10095_),
    .B1(_10097_),
    .B2(_10042_),
    .ZN(_10098_));
 OAI21_X1 _33911_ (.A(_10092_),
    .B1(_10094_),
    .B2(_10098_),
    .ZN(_10099_));
 AOI21_X1 _33912_ (.A(_10087_),
    .B1(_10091_),
    .B2(_10099_),
    .ZN(_10100_));
 INV_X1 _33913_ (.A(_20303_),
    .ZN(_10101_));
 OAI21_X1 _33914_ (.A(_10078_),
    .B1(_10100_),
    .B2(_10101_),
    .ZN(_10102_));
 AOI21_X1 _33915_ (.A(_20300_),
    .B1(_10077_),
    .B2(_10102_),
    .ZN(_10103_));
 OAI21_X2 _33916_ (.A(_10075_),
    .B1(_10076_),
    .B2(_10103_),
    .ZN(_10104_));
 AOI21_X4 _33917_ (.A(_20296_),
    .B1(_20297_),
    .B2(_10104_),
    .ZN(_10105_));
 AND3_X1 _33918_ (.A1(_10093_),
    .A2(_10042_),
    .A3(_10051_),
    .ZN(_10106_));
 AOI21_X2 _33919_ (.A(_10099_),
    .B1(_10106_),
    .B2(_10056_),
    .ZN(_10107_));
 INV_X1 _33920_ (.A(_10107_),
    .ZN(_10108_));
 AOI21_X2 _33921_ (.A(_10087_),
    .B1(_10091_),
    .B2(_10108_),
    .ZN(_10109_));
 XNOR2_X2 _33922_ (.A(_20303_),
    .B(_10109_),
    .ZN(_10110_));
 INV_X1 _33923_ (.A(_20308_),
    .ZN(_10111_));
 INV_X1 _33924_ (.A(_10082_),
    .ZN(_10112_));
 AOI21_X1 _33925_ (.A(_20310_),
    .B1(_10089_),
    .B2(_20312_),
    .ZN(_10113_));
 NAND2_X1 _33926_ (.A1(_10089_),
    .A2(_10093_),
    .ZN(_10114_));
 AOI21_X1 _33927_ (.A(_10095_),
    .B1(_10042_),
    .B2(_20316_),
    .ZN(_10115_));
 OAI21_X1 _33928_ (.A(_10113_),
    .B1(_10114_),
    .B2(_10115_),
    .ZN(_10116_));
 NAND2_X1 _33929_ (.A1(_10042_),
    .A2(_20317_),
    .ZN(_10117_));
 NOR2_X1 _33930_ (.A1(_10114_),
    .A2(_10117_),
    .ZN(_10118_));
 NAND4_X1 _33931_ (.A1(_10013_),
    .A2(_10015_),
    .A3(_20323_),
    .A4(_10031_),
    .ZN(_10119_));
 INV_X1 _33932_ (.A(_10021_),
    .ZN(_10120_));
 AOI21_X1 _33933_ (.A(_20330_),
    .B1(_20332_),
    .B2(_20331_),
    .ZN(_10121_));
 OAI21_X1 _33934_ (.A(_10120_),
    .B1(_10121_),
    .B2(_10061_),
    .ZN(_10122_));
 AOI21_X1 _33935_ (.A(_20326_),
    .B1(_10122_),
    .B2(_10027_),
    .ZN(_10123_));
 OAI221_X1 _33936_ (.A(_10014_),
    .B1(_10016_),
    .B2(_10018_),
    .C1(_10119_),
    .C2(_10123_),
    .ZN(_10124_));
 AOI21_X1 _33937_ (.A(_10116_),
    .B1(_10118_),
    .B2(_10124_),
    .ZN(_10125_));
 OAI21_X1 _33938_ (.A(_10111_),
    .B1(_10112_),
    .B2(_10125_),
    .ZN(_10126_));
 AOI21_X1 _33939_ (.A(_20306_),
    .B1(_10126_),
    .B2(_10085_),
    .ZN(_10127_));
 OAI21_X1 _33940_ (.A(_10079_),
    .B1(_10081_),
    .B2(_10127_),
    .ZN(_10128_));
 AOI21_X2 _33941_ (.A(_20302_),
    .B1(_10128_),
    .B2(_20303_),
    .ZN(_10129_));
 XNOR2_X2 _33942_ (.A(_10077_),
    .B(_10129_),
    .ZN(_10130_));
 AOI21_X2 _33943_ (.A(_20312_),
    .B1(_10093_),
    .B2(_10095_),
    .ZN(_10131_));
 NAND4_X2 _33944_ (.A1(_10082_),
    .A2(_10089_),
    .A3(_10093_),
    .A4(_10042_),
    .ZN(_10132_));
 OAI221_X2 _33945_ (.A(_10083_),
    .B1(_10090_),
    .B2(_10131_),
    .C1(_10132_),
    .C2(_10059_),
    .ZN(_10133_));
 XNOR2_X2 _33946_ (.A(_10088_),
    .B(_10133_),
    .ZN(_10134_));
 INV_X1 _33947_ (.A(_10134_),
    .ZN(_10135_));
 NOR2_X1 _33948_ (.A1(_10016_),
    .A2(_10117_),
    .ZN(_10136_));
 OAI21_X2 _33949_ (.A(_10043_),
    .B1(_10044_),
    .B2(_10014_),
    .ZN(_10137_));
 AOI221_X2 _33950_ (.A(_10095_),
    .B1(_10039_),
    .B2(_10136_),
    .C1(_10137_),
    .C2(_10042_),
    .ZN(_10138_));
 XNOR2_X2 _33951_ (.A(_10093_),
    .B(_10138_),
    .ZN(_10139_));
 NAND3_X1 _33952_ (.A1(_10035_),
    .A2(_20349_),
    .A3(_10139_),
    .ZN(_10140_));
 NOR3_X1 _33953_ (.A1(_10034_),
    .A2(_10114_),
    .A3(_10117_),
    .ZN(_10141_));
 NOR2_X1 _33954_ (.A1(_10116_),
    .A2(_10141_),
    .ZN(_10142_));
 XNOR2_X2 _33955_ (.A(_10112_),
    .B(_10142_),
    .ZN(_10143_));
 XOR2_X2 _33956_ (.A(_10089_),
    .B(_10107_),
    .Z(_10144_));
 OR3_X1 _33957_ (.A1(_10140_),
    .A2(_10143_),
    .A3(_10144_),
    .ZN(_10145_));
 OAI21_X1 _33958_ (.A(_10111_),
    .B1(_10112_),
    .B2(_10113_),
    .ZN(_10146_));
 AOI21_X1 _33959_ (.A(_20306_),
    .B1(_10146_),
    .B2(_10085_),
    .ZN(_10147_));
 NAND4_X1 _33960_ (.A1(_10085_),
    .A2(_10082_),
    .A3(_10089_),
    .A4(_10093_),
    .ZN(_10148_));
 OAI21_X1 _33961_ (.A(_10147_),
    .B1(_10148_),
    .B2(_10138_),
    .ZN(_10149_));
 XNOR2_X2 _33962_ (.A(_10080_),
    .B(_10149_),
    .ZN(_10150_));
 NOR3_X1 _33963_ (.A1(_10135_),
    .A2(_10145_),
    .A3(_10150_),
    .ZN(_10151_));
 NAND3_X2 _33964_ (.A1(_10110_),
    .A2(_10130_),
    .A3(_10151_),
    .ZN(_10152_));
 AOI21_X1 _33965_ (.A(_10021_),
    .B1(_20330_),
    .B2(_20329_),
    .ZN(_10153_));
 OAI21_X1 _33966_ (.A(_10052_),
    .B1(_10055_),
    .B2(_10153_),
    .ZN(_10154_));
 AOI21_X1 _33967_ (.A(_10048_),
    .B1(_10051_),
    .B2(_10154_),
    .ZN(_10155_));
 OAI221_X1 _33968_ (.A(_10083_),
    .B1(_10090_),
    .B2(_10131_),
    .C1(_10132_),
    .C2(_10155_),
    .ZN(_10156_));
 AOI21_X1 _33969_ (.A(_20306_),
    .B1(_10156_),
    .B2(_10085_),
    .ZN(_10157_));
 INV_X1 _33970_ (.A(_10157_),
    .ZN(_10158_));
 AOI21_X1 _33971_ (.A(_20304_),
    .B1(_10080_),
    .B2(_10158_),
    .ZN(_10159_));
 OAI21_X1 _33972_ (.A(_10078_),
    .B1(_10159_),
    .B2(_10101_),
    .ZN(_10160_));
 AOI21_X2 _33973_ (.A(_20300_),
    .B1(_10077_),
    .B2(_10160_),
    .ZN(_10161_));
 XNOR2_X2 _33974_ (.A(_10076_),
    .B(_10161_),
    .ZN(_10162_));
 AOI21_X1 _33975_ (.A(_20326_),
    .B1(_10021_),
    .B2(_10027_),
    .ZN(_10163_));
 INV_X1 _33976_ (.A(_10163_),
    .ZN(_10164_));
 AOI21_X1 _33977_ (.A(_10017_),
    .B1(_10031_),
    .B2(_10164_),
    .ZN(_10165_));
 OAI21_X1 _33978_ (.A(_10037_),
    .B1(_10165_),
    .B2(_10030_),
    .ZN(_10166_));
 AOI221_X2 _33979_ (.A(_10095_),
    .B1(_10136_),
    .B2(_10166_),
    .C1(_10137_),
    .C2(_10042_),
    .ZN(_10167_));
 OAI21_X1 _33980_ (.A(_10147_),
    .B1(_10148_),
    .B2(_10167_),
    .ZN(_10168_));
 AOI21_X1 _33981_ (.A(_20304_),
    .B1(_10080_),
    .B2(_10168_),
    .ZN(_10169_));
 OAI21_X1 _33982_ (.A(_10078_),
    .B1(_10169_),
    .B2(_10101_),
    .ZN(_10170_));
 AOI21_X1 _33983_ (.A(_20300_),
    .B1(_10077_),
    .B2(_10170_),
    .ZN(_10171_));
 OAI21_X1 _33984_ (.A(_10075_),
    .B1(_10076_),
    .B2(_10171_),
    .ZN(_10172_));
 XNOR2_X2 _33985_ (.A(_20297_),
    .B(_10172_),
    .ZN(_10173_));
 NOR3_X1 _33986_ (.A1(_10152_),
    .A2(_10162_),
    .A3(_10173_),
    .ZN(_10174_));
 XOR2_X2 _33987_ (.A(_10105_),
    .B(_10174_),
    .Z(_10175_));
 BUF_X1 _33988_ (.A(_10175_),
    .Z(_14483_));
 OR4_X1 _33989_ (.A1(\g_row[3].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_10176_));
 OAI21_X2 _33990_ (.A(_07621_),
    .B1(_10176_),
    .B2(\g_row[3].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_10177_));
 AND4_X1 _33991_ (.A1(\g_row[3].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .A2(\g_row[3].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .A3(\g_row[3].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .A4(\g_row[3].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .ZN(_10178_));
 AOI21_X4 _33992_ (.A(_07625_),
    .B1(_10178_),
    .B2(\g_row[3].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .ZN(_10179_));
 INV_X1 _33993_ (.A(_14482_),
    .ZN(_10180_));
 AOI21_X1 _33994_ (.A(_10177_),
    .B1(_10179_),
    .B2(_10180_),
    .ZN(_00433_));
 INV_X1 _33995_ (.A(_20339_),
    .ZN(_10181_));
 AOI21_X1 _33996_ (.A(_10177_),
    .B1(_10179_),
    .B2(_10181_),
    .ZN(_00434_));
 INV_X1 _33997_ (.A(_14490_),
    .ZN(_10182_));
 AOI21_X1 _33998_ (.A(_10177_),
    .B1(_10179_),
    .B2(_10182_),
    .ZN(_00435_));
 XOR2_X1 _33999_ (.A(_14489_),
    .B(_20348_),
    .Z(_10183_));
 AOI21_X1 _34000_ (.A(_10177_),
    .B1(_10179_),
    .B2(_10183_),
    .ZN(_00436_));
 AOI21_X1 _34001_ (.A(_20343_),
    .B1(_20344_),
    .B2(_20338_),
    .ZN(_10184_));
 INV_X1 _34002_ (.A(_10184_),
    .ZN(_10185_));
 AOI21_X1 _34003_ (.A(_20347_),
    .B1(_10185_),
    .B2(_20348_),
    .ZN(_10186_));
 XNOR2_X1 _34004_ (.A(\g_row[3].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .B(_20345_),
    .ZN(_10187_));
 XNOR2_X1 _34005_ (.A(_07619_),
    .B(_10187_),
    .ZN(_10188_));
 XNOR2_X1 _34006_ (.A(_10186_),
    .B(_10188_),
    .ZN(_10189_));
 AOI21_X1 _34007_ (.A(_10177_),
    .B1(_10179_),
    .B2(_10189_),
    .ZN(_00437_));
 INV_X1 _34008_ (.A(_10177_),
    .ZN(_10190_));
 NAND2_X4 _34009_ (.A1(_10190_),
    .A2(_10179_),
    .ZN(_10191_));
 INV_X1 _34010_ (.A(_10175_),
    .ZN(_14479_));
 NAND2_X1 _34011_ (.A1(_20352_),
    .A2(_14479_),
    .ZN(_10192_));
 NAND3_X1 _34012_ (.A1(_10035_),
    .A2(_10074_),
    .A3(_14483_),
    .ZN(_10193_));
 AOI21_X2 _34013_ (.A(_10191_),
    .B1(_10192_),
    .B2(_10193_),
    .ZN(_00432_));
 XNOR2_X1 _34014_ (.A(_20351_),
    .B(_10139_),
    .ZN(_10194_));
 INV_X1 _34015_ (.A(_20352_),
    .ZN(_10195_));
 MUX2_X1 _34016_ (.A(_10194_),
    .B(_10195_),
    .S(_14483_),
    .Z(_10196_));
 NOR2_X1 _34017_ (.A1(_10191_),
    .A2(_10196_),
    .ZN(_00438_));
 XNOR2_X1 _34018_ (.A(_10140_),
    .B(_10144_),
    .ZN(_10197_));
 MUX2_X1 _34019_ (.A(_10197_),
    .B(_10194_),
    .S(_14483_),
    .Z(_10198_));
 NOR2_X1 _34020_ (.A1(_10191_),
    .A2(_10198_),
    .ZN(_00439_));
 INV_X1 _34021_ (.A(_10143_),
    .ZN(_10199_));
 INV_X1 _34022_ (.A(_10144_),
    .ZN(_10200_));
 AND3_X1 _34023_ (.A1(_20351_),
    .A2(_10139_),
    .A3(_10200_),
    .ZN(_10201_));
 XNOR2_X1 _34024_ (.A(_10199_),
    .B(_10201_),
    .ZN(_10202_));
 MUX2_X1 _34025_ (.A(_10202_),
    .B(_10197_),
    .S(_14483_),
    .Z(_10203_));
 NOR2_X1 _34026_ (.A1(_10191_),
    .A2(_10203_),
    .ZN(_00440_));
 XNOR2_X1 _34027_ (.A(_10135_),
    .B(_10145_),
    .ZN(_10204_));
 MUX2_X1 _34028_ (.A(_10204_),
    .B(_10202_),
    .S(_14483_),
    .Z(_10205_));
 NOR2_X1 _34029_ (.A1(_10191_),
    .A2(_10205_),
    .ZN(_00441_));
 AND3_X1 _34030_ (.A1(_10134_),
    .A2(_10199_),
    .A3(_10201_),
    .ZN(_10206_));
 XOR2_X1 _34031_ (.A(_10150_),
    .B(_10206_),
    .Z(_10207_));
 MUX2_X1 _34032_ (.A(_10207_),
    .B(_10204_),
    .S(_14483_),
    .Z(_10208_));
 NOR2_X1 _34033_ (.A1(_10191_),
    .A2(_10208_),
    .ZN(_00442_));
 XNOR2_X1 _34034_ (.A(_10110_),
    .B(_10151_),
    .ZN(_10209_));
 MUX2_X1 _34035_ (.A(_10209_),
    .B(_10207_),
    .S(_14483_),
    .Z(_10210_));
 NOR2_X1 _34036_ (.A1(_10191_),
    .A2(_10210_),
    .ZN(_00443_));
 NAND2_X1 _34037_ (.A1(_10110_),
    .A2(_10206_),
    .ZN(_10211_));
 NOR2_X1 _34038_ (.A1(_10150_),
    .A2(_10211_),
    .ZN(_10212_));
 XNOR2_X1 _34039_ (.A(_10130_),
    .B(_10212_),
    .ZN(_10213_));
 MUX2_X1 _34040_ (.A(_10213_),
    .B(_10209_),
    .S(_14483_),
    .Z(_10214_));
 NOR2_X1 _34041_ (.A1(_10191_),
    .A2(_10214_),
    .ZN(_00444_));
 XNOR2_X1 _34042_ (.A(_10152_),
    .B(_10162_),
    .ZN(_10215_));
 MUX2_X1 _34043_ (.A(_10215_),
    .B(_10213_),
    .S(_10175_),
    .Z(_10216_));
 NOR2_X1 _34044_ (.A1(_10191_),
    .A2(_10216_),
    .ZN(_00445_));
 AND2_X1 _34045_ (.A1(_10130_),
    .A2(_10212_),
    .ZN(_10217_));
 OR3_X1 _34046_ (.A1(_10173_),
    .A2(_14483_),
    .A3(_10217_),
    .ZN(_10218_));
 NAND2_X1 _34047_ (.A1(_10173_),
    .A2(_10217_),
    .ZN(_10219_));
 NAND2_X1 _34048_ (.A1(_14479_),
    .A2(_10219_),
    .ZN(_10220_));
 OAI21_X1 _34049_ (.A(_10220_),
    .B1(_14479_),
    .B2(_10152_),
    .ZN(_10221_));
 MUX2_X1 _34050_ (.A(_10173_),
    .B(_10152_),
    .S(_10105_),
    .Z(_10222_));
 MUX2_X1 _34051_ (.A(_10221_),
    .B(_10222_),
    .S(_10162_),
    .Z(_10223_));
 AOI21_X1 _34052_ (.A(_10191_),
    .B1(_10218_),
    .B2(_10223_),
    .ZN(_00446_));
 BUF_X2 _34053_ (.A(\g_reduce0[0].adder.a[12] ),
    .Z(_10224_));
 BUF_X2 _34054_ (.A(\g_reduce0[0].adder.a[14] ),
    .Z(_10225_));
 OR2_X2 _34055_ (.A1(\g_reduce0[0].adder.a[10] ),
    .A2(\g_reduce0[0].adder.a[13] ),
    .ZN(_10226_));
 NOR4_X4 _34056_ (.A1(\g_reduce0[0].adder.a[11] ),
    .A2(_10224_),
    .A3(_10225_),
    .A4(_10226_),
    .ZN(_10227_));
 BUF_X2 _34057_ (.A(\g_reduce0[0].adder.b[14] ),
    .Z(_10228_));
 OR2_X1 _34058_ (.A1(\g_reduce0[0].adder.b[10] ),
    .A2(\g_reduce0[0].adder.b[13] ),
    .ZN(_10229_));
 OR4_X1 _34059_ (.A1(\g_reduce0[0].adder.b[11] ),
    .A2(\g_reduce0[0].adder.b[12] ),
    .A3(_10228_),
    .A4(_10229_),
    .ZN(_10230_));
 BUF_X4 _34060_ (.A(_10230_),
    .Z(_10231_));
 BUF_X2 _34061_ (.A(_20394_),
    .Z(_10232_));
 BUF_X1 _34062_ (.A(_20361_),
    .Z(_10233_));
 BUF_X4 _34063_ (.A(_20355_),
    .Z(_10234_));
 BUF_X2 _34064_ (.A(_20358_),
    .Z(_10235_));
 AND2_X1 _34065_ (.A1(_10234_),
    .A2(_10235_),
    .ZN(_10236_));
 BUF_X4 _34066_ (.A(_10236_),
    .Z(_10237_));
 NAND4_X4 _34067_ (.A1(_20400_),
    .A2(_10232_),
    .A3(_10233_),
    .A4(_10237_),
    .ZN(_10238_));
 AND4_X2 _34068_ (.A1(_20376_),
    .A2(_20379_),
    .A3(_20382_),
    .A4(_20385_),
    .ZN(_10239_));
 AND4_X2 _34069_ (.A1(_20364_),
    .A2(_20367_),
    .A3(_20370_),
    .A4(_20373_),
    .ZN(_10240_));
 NAND4_X4 _34070_ (.A1(_20388_),
    .A2(_20391_),
    .A3(_10239_),
    .A4(_10240_),
    .ZN(_10241_));
 AOI21_X2 _34071_ (.A(_20363_),
    .B1(_20366_),
    .B2(_20364_),
    .ZN(_10242_));
 NAND2_X1 _34072_ (.A1(_20364_),
    .A2(_20367_),
    .ZN(_10243_));
 AOI21_X2 _34073_ (.A(_20369_),
    .B1(_20370_),
    .B2(_20372_),
    .ZN(_10244_));
 OAI21_X4 _34074_ (.A(_10242_),
    .B1(_10243_),
    .B2(_10244_),
    .ZN(_10245_));
 AOI21_X4 _34075_ (.A(_10238_),
    .B1(_10241_),
    .B2(_10245_),
    .ZN(_10246_));
 NAND3_X2 _34076_ (.A1(_20388_),
    .A2(_20391_),
    .A3(_10239_),
    .ZN(_10247_));
 NAND2_X4 _34077_ (.A1(_10240_),
    .A2(_10247_),
    .ZN(_10248_));
 INV_X1 _34078_ (.A(_20387_),
    .ZN(_10249_));
 INV_X1 _34079_ (.A(_20388_),
    .ZN(_10250_));
 OAI21_X1 _34080_ (.A(_10249_),
    .B1(_20390_),
    .B2(_10250_),
    .ZN(_10251_));
 INV_X1 _34081_ (.A(_20378_),
    .ZN(_10252_));
 AOI21_X1 _34082_ (.A(_20381_),
    .B1(_20382_),
    .B2(_20384_),
    .ZN(_10253_));
 INV_X1 _34083_ (.A(_20379_),
    .ZN(_10254_));
 OAI21_X1 _34084_ (.A(_10252_),
    .B1(_10253_),
    .B2(_10254_),
    .ZN(_10255_));
 AOI221_X2 _34085_ (.A(_20375_),
    .B1(_10239_),
    .B2(_10251_),
    .C1(_10255_),
    .C2(_20376_),
    .ZN(_10256_));
 OAI21_X4 _34086_ (.A(_10246_),
    .B1(_10248_),
    .B2(_10256_),
    .ZN(_10257_));
 BUF_X2 _34087_ (.A(_20399_),
    .Z(_10258_));
 INV_X2 _34088_ (.A(_10258_),
    .ZN(_10259_));
 INV_X1 _34089_ (.A(_20360_),
    .ZN(_10260_));
 INV_X1 _34090_ (.A(_10233_),
    .ZN(_10261_));
 OAI21_X1 _34091_ (.A(_10260_),
    .B1(_20393_),
    .B2(_10261_),
    .ZN(_10262_));
 AOI221_X1 _34092_ (.A(_20354_),
    .B1(_10237_),
    .B2(_10262_),
    .C1(_20357_),
    .C2(_10234_),
    .ZN(_10263_));
 BUF_X1 _34093_ (.A(_10263_),
    .Z(_10264_));
 BUF_X4 _34094_ (.A(_20400_),
    .Z(_10265_));
 INV_X2 _34095_ (.A(_10265_),
    .ZN(_10266_));
 OAI211_X4 _34096_ (.A(_10259_),
    .B(_10238_),
    .C1(_10264_),
    .C2(_10266_),
    .ZN(_10267_));
 NAND2_X1 _34097_ (.A1(_10257_),
    .A2(_10267_),
    .ZN(_10268_));
 AOI21_X1 _34098_ (.A(net344),
    .B1(_10231_),
    .B2(_10268_),
    .ZN(_10269_));
 MUX2_X1 _34099_ (.A(\g_reduce0[0].adder.b[15] ),
    .B(\g_reduce0[0].adder.a[15] ),
    .S(_10269_),
    .Z(_00006_));
 BUF_X1 _34100_ (.A(_20392_),
    .Z(_10270_));
 AND2_X1 _34101_ (.A1(_10257_),
    .A2(_10267_),
    .ZN(_10271_));
 BUF_X2 _34102_ (.A(_10271_),
    .Z(_10272_));
 BUF_X4 _34103_ (.A(_10272_),
    .Z(_10273_));
 MUX2_X2 _34104_ (.A(_00450_),
    .B(_10270_),
    .S(_10273_),
    .Z(_20478_));
 MUX2_X2 _34105_ (.A(_20359_),
    .B(_00453_),
    .S(_10273_),
    .Z(_14500_));
 NOR2_X1 _34106_ (.A1(_10245_),
    .A2(_10240_),
    .ZN(_10274_));
 INV_X1 _34107_ (.A(_10245_),
    .ZN(_10275_));
 AOI21_X4 _34108_ (.A(_10274_),
    .B1(_10256_),
    .B2(_10275_),
    .ZN(_10276_));
 AND4_X1 _34109_ (.A1(_20400_),
    .A2(_10232_),
    .A3(_10233_),
    .A4(_10237_),
    .ZN(_10277_));
 BUF_X4 _34110_ (.A(_10277_),
    .Z(_10278_));
 NOR2_X1 _34111_ (.A1(\g_reduce0[0].adder.b[12] ),
    .A2(_00458_),
    .ZN(_10279_));
 AND3_X1 _34112_ (.A1(_10278_),
    .A2(_10241_),
    .A3(_10279_),
    .ZN(_10280_));
 AND2_X4 _34113_ (.A1(_10276_),
    .A2(_10280_),
    .ZN(_10281_));
 NOR2_X2 _34114_ (.A1(_10224_),
    .A2(_20356_),
    .ZN(_10282_));
 OAI211_X4 _34115_ (.A(_10246_),
    .B(_10282_),
    .C1(_10256_),
    .C2(_10248_),
    .ZN(_10283_));
 AND2_X1 _34116_ (.A1(_10238_),
    .A2(_10282_),
    .ZN(_10284_));
 OAI211_X2 _34117_ (.A(_10259_),
    .B(_10284_),
    .C1(_10264_),
    .C2(_10266_),
    .ZN(_10285_));
 NAND2_X1 _34118_ (.A1(_10238_),
    .A2(_10279_),
    .ZN(_10286_));
 AOI21_X2 _34119_ (.A(_20354_),
    .B1(_20357_),
    .B2(_10234_),
    .ZN(_10287_));
 INV_X1 _34120_ (.A(_20393_),
    .ZN(_10288_));
 AOI21_X2 _34121_ (.A(_20360_),
    .B1(_10288_),
    .B2(_10233_),
    .ZN(_10289_));
 INV_X1 _34122_ (.A(_10237_),
    .ZN(_10290_));
 OAI21_X4 _34123_ (.A(_10287_),
    .B1(_10289_),
    .B2(_10290_),
    .ZN(_10291_));
 AOI21_X4 _34124_ (.A(_10258_),
    .B1(_10291_),
    .B2(_10265_),
    .ZN(_10292_));
 OAI211_X4 _34125_ (.A(_10283_),
    .B(_10285_),
    .C1(_10286_),
    .C2(_10292_),
    .ZN(_10293_));
 OR2_X2 _34126_ (.A1(\g_reduce0[0].adder.a[11] ),
    .A2(_20359_),
    .ZN(_10294_));
 NOR2_X1 _34127_ (.A1(_10278_),
    .A2(_10294_),
    .ZN(_10295_));
 OAI211_X2 _34128_ (.A(_10259_),
    .B(_10295_),
    .C1(_10264_),
    .C2(_10266_),
    .ZN(_10296_));
 NOR2_X1 _34129_ (.A1(\g_reduce0[0].adder.b[11] ),
    .A2(_00453_),
    .ZN(_10297_));
 NAND3_X1 _34130_ (.A1(_10278_),
    .A2(_10241_),
    .A3(_10297_),
    .ZN(_10298_));
 AND3_X1 _34131_ (.A1(_20376_),
    .A2(_10255_),
    .A3(_10240_),
    .ZN(_10299_));
 INV_X1 _34132_ (.A(_20375_),
    .ZN(_10300_));
 INV_X1 _34133_ (.A(_10239_),
    .ZN(_10301_));
 INV_X1 _34134_ (.A(_20390_),
    .ZN(_10302_));
 AOI21_X1 _34135_ (.A(_20387_),
    .B1(_10302_),
    .B2(_20388_),
    .ZN(_10303_));
 OAI21_X1 _34136_ (.A(_10300_),
    .B1(_10301_),
    .B2(_10303_),
    .ZN(_10304_));
 AOI211_X2 _34137_ (.A(_10245_),
    .B(_10299_),
    .C1(_10240_),
    .C2(_10304_),
    .ZN(_10305_));
 NAND2_X1 _34138_ (.A1(_10238_),
    .A2(_10297_),
    .ZN(_10306_));
 OAI221_X2 _34139_ (.A(_10296_),
    .B1(_10298_),
    .B2(_10305_),
    .C1(_10292_),
    .C2(_10306_),
    .ZN(_10307_));
 INV_X1 _34140_ (.A(_20396_),
    .ZN(_10308_));
 AOI211_X2 _34141_ (.A(_10238_),
    .B(_10294_),
    .C1(_10241_),
    .C2(_10245_),
    .ZN(_10309_));
 OAI21_X4 _34142_ (.A(_10309_),
    .B1(_10248_),
    .B2(_10256_),
    .ZN(_10310_));
 NAND2_X4 _34143_ (.A1(_10308_),
    .A2(_10310_),
    .ZN(_10311_));
 NOR4_X4 _34144_ (.A1(_10281_),
    .A2(_10293_),
    .A3(_10307_),
    .A4(_10311_),
    .ZN(_10312_));
 NOR3_X1 _34145_ (.A1(\g_reduce0[0].adder.a[13] ),
    .A2(_20353_),
    .A3(_10278_),
    .ZN(_10313_));
 OAI211_X2 _34146_ (.A(_10259_),
    .B(_10313_),
    .C1(_10264_),
    .C2(_10266_),
    .ZN(_10314_));
 NOR2_X1 _34147_ (.A1(\g_reduce0[0].adder.b[13] ),
    .A2(_00461_),
    .ZN(_10315_));
 NAND3_X1 _34148_ (.A1(_10278_),
    .A2(_10241_),
    .A3(_10315_),
    .ZN(_10316_));
 NAND2_X1 _34149_ (.A1(_10238_),
    .A2(_10315_),
    .ZN(_10317_));
 OAI221_X2 _34150_ (.A(_10314_),
    .B1(_10316_),
    .B2(_10305_),
    .C1(_10292_),
    .C2(_10317_),
    .ZN(_10318_));
 NOR3_X4 _34151_ (.A1(\g_reduce0[0].adder.a[13] ),
    .A2(_20353_),
    .A3(_10257_),
    .ZN(_10319_));
 NOR3_X2 _34152_ (.A1(_10265_),
    .A2(_10318_),
    .A3(_10319_),
    .ZN(_10320_));
 NOR2_X1 _34153_ (.A1(_10265_),
    .A2(_10235_),
    .ZN(_10321_));
 NOR4_X4 _34154_ (.A1(_10318_),
    .A2(_10319_),
    .A3(_10281_),
    .A4(_10293_),
    .ZN(_10322_));
 AOI22_X4 _34155_ (.A1(_10312_),
    .A2(_10320_),
    .B1(_10321_),
    .B2(_10322_),
    .ZN(_10323_));
 OAI21_X2 _34156_ (.A(_10265_),
    .B1(_10318_),
    .B2(_10319_),
    .ZN(_10324_));
 OR4_X2 _34157_ (.A1(_10265_),
    .A2(_10234_),
    .A3(_10318_),
    .A4(_10319_),
    .ZN(_10325_));
 INV_X1 _34158_ (.A(_10234_),
    .ZN(_10326_));
 NOR2_X1 _34159_ (.A1(_10266_),
    .A2(_10326_),
    .ZN(_10327_));
 OAI21_X2 _34160_ (.A(_10327_),
    .B1(_10293_),
    .B2(_10281_),
    .ZN(_10328_));
 AND2_X1 _34161_ (.A1(_10235_),
    .A2(_10327_),
    .ZN(_10329_));
 OAI21_X2 _34162_ (.A(_10329_),
    .B1(_10311_),
    .B2(_10307_),
    .ZN(_10330_));
 AND4_X2 _34163_ (.A1(_10324_),
    .A2(_10325_),
    .A3(_10328_),
    .A4(_10330_),
    .ZN(_10331_));
 NAND2_X2 _34164_ (.A1(_10323_),
    .A2(_10331_),
    .ZN(_10332_));
 CLKBUF_X3 _34165_ (.A(_10232_),
    .Z(_10333_));
 MUX2_X1 _34166_ (.A(_00457_),
    .B(_20371_),
    .S(_10273_),
    .Z(_10334_));
 MUX2_X1 _34167_ (.A(_00455_),
    .B(_20377_),
    .S(_10273_),
    .Z(_10335_));
 BUF_X2 _34168_ (.A(_20397_),
    .Z(_10336_));
 INV_X2 _34169_ (.A(_10336_),
    .ZN(_10337_));
 MUX2_X1 _34170_ (.A(_10334_),
    .B(_10335_),
    .S(_10337_),
    .Z(_10338_));
 NAND2_X1 _34171_ (.A1(_10333_),
    .A2(_10338_),
    .ZN(_10339_));
 AND2_X1 _34172_ (.A1(_00454_),
    .A2(_10268_),
    .ZN(_10340_));
 AOI21_X1 _34173_ (.A(_10340_),
    .B1(_10273_),
    .B2(_20374_),
    .ZN(_10341_));
 NAND2_X1 _34174_ (.A1(_10337_),
    .A2(_10341_),
    .ZN(_10342_));
 MUX2_X1 _34175_ (.A(_00456_),
    .B(_20368_),
    .S(_10272_),
    .Z(_10343_));
 OAI21_X1 _34176_ (.A(_10342_),
    .B1(_10343_),
    .B2(_10337_),
    .ZN(_10344_));
 OAI21_X1 _34177_ (.A(_10339_),
    .B1(_10344_),
    .B2(_10333_),
    .ZN(_10345_));
 INV_X1 _34178_ (.A(_00450_),
    .ZN(_10346_));
 AND4_X1 _34179_ (.A1(_10346_),
    .A2(_10270_),
    .A3(_10257_),
    .A4(_10267_),
    .ZN(_10347_));
 OR2_X1 _34180_ (.A1(_10346_),
    .A2(_10270_),
    .ZN(_10348_));
 AOI21_X1 _34181_ (.A(_10348_),
    .B1(_10267_),
    .B2(_10257_),
    .ZN(_10349_));
 NAND2_X1 _34182_ (.A1(_10233_),
    .A2(_10237_),
    .ZN(_10350_));
 NOR3_X1 _34183_ (.A1(_10347_),
    .A2(_10349_),
    .A3(_10350_),
    .ZN(_10351_));
 NAND4_X1 _34184_ (.A1(_10346_),
    .A2(_10270_),
    .A3(_10257_),
    .A4(_10267_),
    .ZN(_10352_));
 NOR2_X1 _34185_ (.A1(_10346_),
    .A2(_10270_),
    .ZN(_10353_));
 NAND2_X1 _34186_ (.A1(_10278_),
    .A2(_10241_),
    .ZN(_10354_));
 OAI221_X2 _34187_ (.A(_10353_),
    .B1(_10292_),
    .B2(_10278_),
    .C1(_10305_),
    .C2(_10354_),
    .ZN(_10355_));
 AOI21_X1 _34188_ (.A(_10234_),
    .B1(_10352_),
    .B2(_10355_),
    .ZN(_10356_));
 NOR2_X2 _34189_ (.A1(_10257_),
    .A2(_10294_),
    .ZN(_10357_));
 NOR4_X4 _34190_ (.A1(_10281_),
    .A2(_10293_),
    .A3(_10307_),
    .A4(_10357_),
    .ZN(_10358_));
 NAND2_X1 _34191_ (.A1(_10238_),
    .A2(_10282_),
    .ZN(_10359_));
 AOI211_X2 _34192_ (.A(_10258_),
    .B(_10359_),
    .C1(_10291_),
    .C2(_10265_),
    .ZN(_10360_));
 AND2_X1 _34193_ (.A1(_10238_),
    .A2(_10279_),
    .ZN(_10361_));
 OAI21_X2 _34194_ (.A(_10259_),
    .B1(_10264_),
    .B2(_10266_),
    .ZN(_10362_));
 AOI221_X2 _34195_ (.A(_10360_),
    .B1(_10361_),
    .B2(_10362_),
    .C1(_10276_),
    .C2(_10280_),
    .ZN(_10363_));
 NAND2_X2 _34196_ (.A1(_10283_),
    .A2(_10363_),
    .ZN(_10364_));
 AOI221_X2 _34197_ (.A(_10351_),
    .B1(_10356_),
    .B2(_10358_),
    .C1(_10234_),
    .C2(_10364_),
    .ZN(_10365_));
 OR2_X1 _34198_ (.A1(_10234_),
    .A2(_10235_),
    .ZN(_10366_));
 NOR3_X1 _34199_ (.A1(_10281_),
    .A2(_10293_),
    .A3(_10366_),
    .ZN(_10367_));
 NOR2_X1 _34200_ (.A1(_10234_),
    .A2(_10233_),
    .ZN(_10368_));
 OR2_X1 _34201_ (.A1(_10278_),
    .A2(_10294_),
    .ZN(_10369_));
 AOI211_X2 _34202_ (.A(_10258_),
    .B(_10369_),
    .C1(_10291_),
    .C2(_10265_),
    .ZN(_10370_));
 AND3_X1 _34203_ (.A1(_10278_),
    .A2(_10241_),
    .A3(_10297_),
    .ZN(_10371_));
 AND2_X1 _34204_ (.A1(_10238_),
    .A2(_10297_),
    .ZN(_10372_));
 AOI221_X2 _34205_ (.A(_10370_),
    .B1(_10371_),
    .B2(_10276_),
    .C1(_10362_),
    .C2(_10372_),
    .ZN(_10373_));
 NAND2_X1 _34206_ (.A1(_10373_),
    .A2(_10310_),
    .ZN(_10374_));
 AOI221_X2 _34207_ (.A(_10367_),
    .B1(_10368_),
    .B2(_10358_),
    .C1(_10237_),
    .C2(_10374_),
    .ZN(_10375_));
 NAND2_X2 _34208_ (.A1(_10365_),
    .A2(_10375_),
    .ZN(_10376_));
 OAI21_X4 _34209_ (.A(_10235_),
    .B1(_10307_),
    .B2(_10311_),
    .ZN(_10377_));
 OR3_X4 _34210_ (.A1(_10235_),
    .A2(_10307_),
    .A3(_10311_),
    .ZN(_10378_));
 AND2_X1 _34211_ (.A1(_10377_),
    .A2(_10378_),
    .ZN(_10379_));
 CLKBUF_X3 _34212_ (.A(_10379_),
    .Z(_10380_));
 NAND2_X1 _34213_ (.A1(_10376_),
    .A2(_10380_),
    .ZN(_10381_));
 INV_X2 _34214_ (.A(_10232_),
    .ZN(_10382_));
 CLKBUF_X3 _34215_ (.A(_10336_),
    .Z(_10383_));
 NAND2_X1 _34216_ (.A1(_10382_),
    .A2(_10383_),
    .ZN(_10384_));
 OAI221_X2 _34217_ (.A(_00459_),
    .B1(_10305_),
    .B2(_10354_),
    .C1(_10292_),
    .C2(_10278_),
    .ZN(_10385_));
 NAND3_X1 _34218_ (.A1(_20362_),
    .A2(_10257_),
    .A3(_10267_),
    .ZN(_10386_));
 NAND3_X1 _34219_ (.A1(_10382_),
    .A2(_10385_),
    .A3(_10386_),
    .ZN(_10387_));
 MUX2_X1 _34220_ (.A(_00460_),
    .B(_20365_),
    .S(_10272_),
    .Z(_10388_));
 OAI21_X1 _34221_ (.A(_10387_),
    .B1(_10388_),
    .B2(_10382_),
    .ZN(_10389_));
 OAI21_X1 _34222_ (.A(_10384_),
    .B1(_10389_),
    .B2(_10383_),
    .ZN(_10390_));
 MUX2_X1 _34223_ (.A(_00448_),
    .B(_20386_),
    .S(_10272_),
    .Z(_10391_));
 NOR2_X1 _34224_ (.A1(_10383_),
    .A2(_10391_),
    .ZN(_10392_));
 AND2_X1 _34225_ (.A1(_00451_),
    .A2(_10268_),
    .ZN(_10393_));
 BUF_X4 _34226_ (.A(_10273_),
    .Z(_10394_));
 AOI21_X1 _34227_ (.A(_10393_),
    .B1(_10394_),
    .B2(_20380_),
    .ZN(_10395_));
 AOI21_X1 _34228_ (.A(_10392_),
    .B1(_10395_),
    .B2(_10383_),
    .ZN(_10396_));
 MUX2_X1 _34229_ (.A(_00452_),
    .B(_20383_),
    .S(_10272_),
    .Z(_10397_));
 MUX2_X1 _34230_ (.A(_20389_),
    .B(_00449_),
    .S(_10272_),
    .Z(_10398_));
 MUX2_X1 _34231_ (.A(_10397_),
    .B(_10398_),
    .S(_10337_),
    .Z(_10399_));
 MUX2_X1 _34232_ (.A(_10396_),
    .B(_10399_),
    .S(_10333_),
    .Z(_10400_));
 MUX2_X1 _34233_ (.A(_10390_),
    .B(_10400_),
    .S(_10376_),
    .Z(_10401_));
 OAI22_X1 _34234_ (.A1(_10345_),
    .A2(_10381_),
    .B1(_10401_),
    .B2(_10380_),
    .ZN(_10402_));
 NAND2_X1 _34235_ (.A1(_10332_),
    .A2(_10402_),
    .ZN(_20464_));
 INV_X1 _34236_ (.A(_20464_),
    .ZN(_20461_));
 MUX2_X1 _34237_ (.A(_10335_),
    .B(_10397_),
    .S(_10337_),
    .Z(_10403_));
 MUX2_X1 _34238_ (.A(_10396_),
    .B(_10403_),
    .S(_10382_),
    .Z(_10404_));
 MUX2_X1 _34239_ (.A(_10334_),
    .B(_10388_),
    .S(_10383_),
    .Z(_10405_));
 NOR2_X1 _34240_ (.A1(_10333_),
    .A2(_10405_),
    .ZN(_10406_));
 AOI21_X1 _34241_ (.A(_10406_),
    .B1(_10344_),
    .B2(_10333_),
    .ZN(_10407_));
 MUX2_X1 _34242_ (.A(_10404_),
    .B(_10407_),
    .S(_10380_),
    .Z(_10408_));
 INV_X1 _34243_ (.A(_10408_),
    .ZN(_10409_));
 NAND2_X1 _34244_ (.A1(_10376_),
    .A2(_10409_),
    .ZN(_10410_));
 NAND2_X4 _34245_ (.A1(_10377_),
    .A2(_10378_),
    .ZN(_10411_));
 NAND2_X1 _34246_ (.A1(_10385_),
    .A2(_10386_),
    .ZN(_10412_));
 AOI21_X2 _34247_ (.A(_10383_),
    .B1(_10412_),
    .B2(_10333_),
    .ZN(_10413_));
 NAND2_X1 _34248_ (.A1(_10411_),
    .A2(_10413_),
    .ZN(_10414_));
 OAI21_X1 _34249_ (.A(_10410_),
    .B1(_10414_),
    .B2(_10376_),
    .ZN(_10415_));
 NAND2_X1 _34250_ (.A1(_10332_),
    .A2(_10415_),
    .ZN(_14497_));
 INV_X1 _34251_ (.A(_14497_),
    .ZN(_14492_));
 OR2_X1 _34252_ (.A1(_10307_),
    .A2(_10311_),
    .ZN(_10416_));
 OR3_X1 _34253_ (.A1(_10265_),
    .A2(_10318_),
    .A3(_10319_),
    .ZN(_10417_));
 OR4_X1 _34254_ (.A1(_10318_),
    .A2(_10319_),
    .A3(_10281_),
    .A4(_10293_),
    .ZN(_10418_));
 OAI33_X1 _34255_ (.A1(_10364_),
    .A2(_10416_),
    .A3(_10417_),
    .B1(_10418_),
    .B2(_10265_),
    .B3(_10235_),
    .ZN(_10419_));
 NAND4_X4 _34256_ (.A1(_10324_),
    .A2(_10325_),
    .A3(_10328_),
    .A4(_10330_),
    .ZN(_10420_));
 OAI21_X1 _34257_ (.A(_10234_),
    .B1(_10281_),
    .B2(_10293_),
    .ZN(_10421_));
 OAI21_X1 _34258_ (.A(_10326_),
    .B1(_10347_),
    .B2(_10349_),
    .ZN(_10422_));
 NAND4_X2 _34259_ (.A1(_10283_),
    .A2(_10363_),
    .A3(_10373_),
    .A4(_10310_),
    .ZN(_10423_));
 NAND2_X1 _34260_ (.A1(_10352_),
    .A2(_10355_),
    .ZN(_10424_));
 OAI221_X2 _34261_ (.A(_10421_),
    .B1(_10422_),
    .B2(_10423_),
    .C1(_10424_),
    .C2(_10350_),
    .ZN(_10425_));
 OAI21_X1 _34262_ (.A(_10237_),
    .B1(_10307_),
    .B2(_10357_),
    .ZN(_10426_));
 NAND2_X1 _34263_ (.A1(_10326_),
    .A2(_10261_),
    .ZN(_10427_));
 OAI221_X2 _34264_ (.A(_10426_),
    .B1(_10427_),
    .B2(_10423_),
    .C1(_10364_),
    .C2(_10366_),
    .ZN(_10428_));
 OAI22_X4 _34265_ (.A1(net343),
    .A2(_10420_),
    .B1(_10425_),
    .B2(_10428_),
    .ZN(_10429_));
 BUF_X4 _34266_ (.A(_10429_),
    .Z(_10430_));
 NOR2_X1 _34267_ (.A1(_10380_),
    .A2(_10430_),
    .ZN(_10431_));
 NAND2_X1 _34268_ (.A1(_10413_),
    .A2(_10431_),
    .ZN(_20416_));
 INV_X1 _34269_ (.A(_20416_),
    .ZN(_20420_));
 OR3_X1 _34270_ (.A1(_10380_),
    .A2(_10390_),
    .A3(_10430_),
    .ZN(_20410_));
 INV_X1 _34271_ (.A(_20410_),
    .ZN(_20413_));
 NAND2_X1 _34272_ (.A1(_10232_),
    .A2(_10336_),
    .ZN(_10432_));
 AOI21_X1 _34273_ (.A(_10432_),
    .B1(_10386_),
    .B2(_10385_),
    .ZN(_10433_));
 NOR2_X2 _34274_ (.A1(_10382_),
    .A2(_10336_),
    .ZN(_10434_));
 NOR2_X1 _34275_ (.A1(_10333_),
    .A2(_10383_),
    .ZN(_10435_));
 AOI221_X2 _34276_ (.A(_10433_),
    .B1(_10434_),
    .B2(_10343_),
    .C1(_10435_),
    .C2(_10388_),
    .ZN(_10436_));
 NAND2_X1 _34277_ (.A1(_10431_),
    .A2(_10436_),
    .ZN(_20444_));
 INV_X1 _34278_ (.A(_20444_),
    .ZN(_20448_));
 AOI22_X4 _34279_ (.A1(_10323_),
    .A2(_10331_),
    .B1(_10365_),
    .B2(_10375_),
    .ZN(_10437_));
 NAND2_X1 _34280_ (.A1(_10383_),
    .A2(_10389_),
    .ZN(_10438_));
 MUX2_X1 _34281_ (.A(_10343_),
    .B(_10334_),
    .S(_10333_),
    .Z(_10439_));
 OAI21_X1 _34282_ (.A(_10438_),
    .B1(_10439_),
    .B2(_10383_),
    .ZN(_10440_));
 MUX2_X1 _34283_ (.A(_10434_),
    .B(_10440_),
    .S(_10411_),
    .Z(_10441_));
 NAND2_X1 _34284_ (.A1(_10437_),
    .A2(_10441_),
    .ZN(_20424_));
 INV_X1 _34285_ (.A(_20424_),
    .ZN(_20427_));
 NAND2_X1 _34286_ (.A1(_10380_),
    .A2(_10413_),
    .ZN(_10442_));
 OAI21_X1 _34287_ (.A(_10442_),
    .B1(_10407_),
    .B2(_10380_),
    .ZN(_10443_));
 AND2_X1 _34288_ (.A1(_10437_),
    .A2(_10443_),
    .ZN(_20430_));
 INV_X1 _34289_ (.A(_20430_),
    .ZN(_20434_));
 MUX2_X1 _34290_ (.A(_10345_),
    .B(_10390_),
    .S(_10380_),
    .Z(_10444_));
 NOR2_X1 _34291_ (.A1(_10430_),
    .A2(_10444_),
    .ZN(_20438_));
 INV_X1 _34292_ (.A(_20438_),
    .ZN(_20441_));
 NAND2_X1 _34293_ (.A1(_10383_),
    .A2(_00457_),
    .ZN(_10445_));
 NAND2_X1 _34294_ (.A1(_10337_),
    .A2(_00455_),
    .ZN(_10446_));
 NAND3_X1 _34295_ (.A1(_10382_),
    .A2(_10445_),
    .A3(_10446_),
    .ZN(_10447_));
 MUX2_X1 _34296_ (.A(_00451_),
    .B(_00454_),
    .S(_10336_),
    .Z(_10448_));
 OAI21_X1 _34297_ (.A(_10447_),
    .B1(_10448_),
    .B2(_10382_),
    .ZN(_10449_));
 AOI21_X1 _34298_ (.A(_10449_),
    .B1(_10267_),
    .B2(_10257_),
    .ZN(_10450_));
 MUX2_X1 _34299_ (.A(_20377_),
    .B(_20371_),
    .S(_10336_),
    .Z(_10451_));
 MUX2_X1 _34300_ (.A(_20380_),
    .B(_20374_),
    .S(_10336_),
    .Z(_10452_));
 MUX2_X1 _34301_ (.A(_10451_),
    .B(_10452_),
    .S(_10333_),
    .Z(_10453_));
 AOI21_X2 _34302_ (.A(_10450_),
    .B1(_10453_),
    .B2(_10273_),
    .ZN(_10454_));
 MUX2_X1 _34303_ (.A(_10436_),
    .B(_10454_),
    .S(_10411_),
    .Z(_10455_));
 AND2_X1 _34304_ (.A1(_10437_),
    .A2(_10455_),
    .ZN(_20454_));
 INV_X1 _34305_ (.A(_20454_),
    .ZN(_20458_));
 NAND2_X1 _34306_ (.A1(_10333_),
    .A2(_10337_),
    .ZN(_10456_));
 AOI21_X4 _34307_ (.A(_10456_),
    .B1(_10378_),
    .B2(_10377_),
    .ZN(_10457_));
 MUX2_X1 _34308_ (.A(_10341_),
    .B(_10395_),
    .S(_10337_),
    .Z(_10458_));
 NAND2_X1 _34309_ (.A1(_10382_),
    .A2(_10458_),
    .ZN(_10459_));
 OAI21_X1 _34310_ (.A(_10459_),
    .B1(_10403_),
    .B2(_10382_),
    .ZN(_10460_));
 MUX2_X1 _34311_ (.A(_10440_),
    .B(_10460_),
    .S(_10411_),
    .Z(_10461_));
 MUX2_X1 _34312_ (.A(_10457_),
    .B(_10461_),
    .S(_10376_),
    .Z(_10462_));
 NAND2_X1 _34313_ (.A1(_10332_),
    .A2(_10462_),
    .ZN(_20451_));
 INV_X1 _34314_ (.A(_20451_),
    .ZN(_20405_));
 NAND2_X4 _34315_ (.A1(_10411_),
    .A2(_10434_),
    .ZN(_10463_));
 XNOR2_X2 _34316_ (.A(\g_reduce0[0].adder.b[15] ),
    .B(\g_reduce0[0].adder.a[15] ),
    .ZN(_10464_));
 CLKBUF_X3 _34317_ (.A(_10464_),
    .Z(_10465_));
 INV_X1 _34318_ (.A(_20411_),
    .ZN(_10466_));
 INV_X1 _34319_ (.A(_20446_),
    .ZN(_10467_));
 INV_X1 _34320_ (.A(_20425_),
    .ZN(_10468_));
 BUF_X1 _34321_ (.A(_20447_),
    .Z(_10469_));
 INV_X1 _34322_ (.A(_10469_),
    .ZN(_10470_));
 OAI21_X2 _34323_ (.A(_10467_),
    .B1(_10468_),
    .B2(_10470_),
    .ZN(_10471_));
 INV_X1 _34324_ (.A(_20435_),
    .ZN(_10472_));
 BUF_X2 _34325_ (.A(_20433_),
    .Z(_10473_));
 BUF_X2 _34326_ (.A(_20440_),
    .Z(_10474_));
 NOR2_X2 _34327_ (.A1(_20435_),
    .A2(_20442_),
    .ZN(_10475_));
 NOR3_X2 _34328_ (.A1(_20435_),
    .A2(_20442_),
    .A3(_20459_),
    .ZN(_10476_));
 INV_X1 _34329_ (.A(_20457_),
    .ZN(_10477_));
 AND2_X1 _34330_ (.A1(_14496_),
    .A2(_20404_),
    .ZN(_10478_));
 OR2_X1 _34331_ (.A1(_20403_),
    .A2(_20452_),
    .ZN(_10479_));
 BUF_X1 _34332_ (.A(_20453_),
    .Z(_10480_));
 OAI221_X2 _34333_ (.A(_10477_),
    .B1(_10478_),
    .B2(_10479_),
    .C1(_10480_),
    .C2(_20452_),
    .ZN(_10481_));
 AOI222_X2 _34334_ (.A1(_10472_),
    .A2(_10473_),
    .B1(_10474_),
    .B2(_10475_),
    .C1(_10476_),
    .C2(_10481_),
    .ZN(_10482_));
 INV_X2 _34335_ (.A(_20426_),
    .ZN(_10483_));
 NOR2_X2 _34336_ (.A1(_10483_),
    .A2(_10470_),
    .ZN(_10484_));
 AOI21_X1 _34337_ (.A(_10471_),
    .B1(_10482_),
    .B2(_10484_),
    .ZN(_10485_));
 INV_X2 _34338_ (.A(_20412_),
    .ZN(_10486_));
 OAI21_X1 _34339_ (.A(_10466_),
    .B1(_10485_),
    .B2(_10486_),
    .ZN(_10487_));
 BUF_X2 _34340_ (.A(_20419_),
    .Z(_10488_));
 AOI21_X1 _34341_ (.A(_20418_),
    .B1(_10487_),
    .B2(_10488_),
    .ZN(_10489_));
 OR2_X2 _34342_ (.A1(_10465_),
    .A2(_10489_),
    .ZN(_10490_));
 XOR2_X2 _34343_ (.A(\g_reduce0[0].adder.b[15] ),
    .B(\g_reduce0[0].adder.a[15] ),
    .Z(_10491_));
 BUF_X4 _34344_ (.A(_10491_),
    .Z(_10492_));
 AOI21_X1 _34345_ (.A(_10488_),
    .B1(_20418_),
    .B2(_10492_),
    .ZN(_10493_));
 OR2_X1 _34346_ (.A1(_20414_),
    .A2(_10492_),
    .ZN(_10494_));
 INV_X1 _34347_ (.A(_20449_),
    .ZN(_10495_));
 OR2_X1 _34348_ (.A1(_20428_),
    .A2(_20432_),
    .ZN(_10496_));
 NOR2_X1 _34349_ (.A1(_20439_),
    .A2(_20456_),
    .ZN(_10497_));
 BUF_X1 _34350_ (.A(_20408_),
    .Z(_10498_));
 AOI21_X1 _34351_ (.A(_20407_),
    .B1(_14494_),
    .B2(_10498_),
    .ZN(_10499_));
 OAI21_X1 _34352_ (.A(_10497_),
    .B1(_10499_),
    .B2(_10477_),
    .ZN(_10500_));
 OR2_X1 _34353_ (.A1(_10474_),
    .A2(_20439_),
    .ZN(_10501_));
 AND2_X1 _34354_ (.A1(_10473_),
    .A2(_10501_),
    .ZN(_10502_));
 AOI21_X1 _34355_ (.A(_10496_),
    .B1(_10500_),
    .B2(_10502_),
    .ZN(_10503_));
 OAI21_X1 _34356_ (.A(_10470_),
    .B1(_20428_),
    .B2(_10483_),
    .ZN(_10504_));
 OAI21_X1 _34357_ (.A(_10495_),
    .B1(_10503_),
    .B2(_10504_),
    .ZN(_10505_));
 AND2_X1 _34358_ (.A1(_10486_),
    .A2(_10505_),
    .ZN(_10506_));
 OAI21_X2 _34359_ (.A(_10493_),
    .B1(_10494_),
    .B2(_10506_),
    .ZN(_10507_));
 NAND2_X2 _34360_ (.A1(_20421_),
    .A2(_10465_),
    .ZN(_10508_));
 NAND2_X1 _34361_ (.A1(_10466_),
    .A2(_10491_),
    .ZN(_10509_));
 NOR2_X1 _34362_ (.A1(_20418_),
    .A2(_10509_),
    .ZN(_10510_));
 AOI21_X1 _34363_ (.A(_20452_),
    .B1(_14498_),
    .B2(_10480_),
    .ZN(_10511_));
 OR2_X1 _34364_ (.A1(_20457_),
    .A2(_10511_),
    .ZN(_10512_));
 AOI222_X1 _34365_ (.A1(_10472_),
    .A2(_10473_),
    .B1(_10474_),
    .B2(_10475_),
    .C1(_10476_),
    .C2(_10512_),
    .ZN(_10513_));
 AOI21_X2 _34366_ (.A(_10471_),
    .B1(_10484_),
    .B2(_10513_),
    .ZN(_10514_));
 OAI21_X2 _34367_ (.A(_10510_),
    .B1(_10514_),
    .B2(_10486_),
    .ZN(_10515_));
 AND3_X2 _34368_ (.A1(_10507_),
    .A2(_10508_),
    .A3(_10515_),
    .ZN(_10516_));
 OR4_X1 _34369_ (.A1(_10430_),
    .A2(_10463_),
    .A3(_10490_),
    .A4(_10516_),
    .ZN(_10517_));
 INV_X1 _34370_ (.A(_20421_),
    .ZN(_10518_));
 OAI21_X1 _34371_ (.A(_20457_),
    .B1(_10498_),
    .B2(_20407_),
    .ZN(_10519_));
 AOI211_X2 _34372_ (.A(_20401_),
    .B(_20407_),
    .C1(_14491_),
    .C2(_20402_),
    .ZN(_10520_));
 OAI21_X1 _34373_ (.A(_10497_),
    .B1(_10519_),
    .B2(_10520_),
    .ZN(_10521_));
 AND3_X1 _34374_ (.A1(_10483_),
    .A2(_10473_),
    .A3(_10501_),
    .ZN(_10522_));
 AOI221_X2 _34375_ (.A(_20428_),
    .B1(_10521_),
    .B2(_10522_),
    .C1(_20432_),
    .C2(_10483_),
    .ZN(_10523_));
 OAI21_X1 _34376_ (.A(_10495_),
    .B1(_10469_),
    .B2(_10523_),
    .ZN(_10524_));
 AOI21_X1 _34377_ (.A(_20414_),
    .B1(_10524_),
    .B2(_10486_),
    .ZN(_10525_));
 OAI21_X2 _34378_ (.A(_10518_),
    .B1(_10488_),
    .B2(_10525_),
    .ZN(_10526_));
 AND2_X1 _34379_ (.A1(_10465_),
    .A2(_10526_),
    .ZN(_10527_));
 NAND3_X4 _34380_ (.A1(_10507_),
    .A2(_10508_),
    .A3(_10515_),
    .ZN(_10528_));
 NOR2_X1 _34381_ (.A1(_10527_),
    .A2(_10528_),
    .ZN(_10529_));
 OAI21_X1 _34382_ (.A(_10529_),
    .B1(_10463_),
    .B2(_10430_),
    .ZN(_10530_));
 NAND2_X1 _34383_ (.A1(_10517_),
    .A2(_10530_),
    .ZN(_10531_));
 AOI211_X2 _34384_ (.A(_10471_),
    .B(_10509_),
    .C1(_10484_),
    .C2(_10482_),
    .ZN(_10532_));
 AOI21_X1 _34385_ (.A(_20412_),
    .B1(_20411_),
    .B2(_10491_),
    .ZN(_10533_));
 NOR2_X1 _34386_ (.A1(_20449_),
    .A2(_10491_),
    .ZN(_10534_));
 OAI21_X1 _34387_ (.A(_10534_),
    .B1(_10523_),
    .B2(_10469_),
    .ZN(_10535_));
 AOI221_X2 _34388_ (.A(_10532_),
    .B1(_10533_),
    .B2(_10535_),
    .C1(_20414_),
    .C2(_10464_),
    .ZN(_10536_));
 XNOR2_X2 _34389_ (.A(_10488_),
    .B(_10536_),
    .ZN(_10537_));
 OR3_X1 _34390_ (.A1(_10483_),
    .A2(_20428_),
    .A3(_10491_),
    .ZN(_10538_));
 OAI21_X1 _34391_ (.A(_10538_),
    .B1(_10464_),
    .B2(_10468_),
    .ZN(_10539_));
 OR2_X1 _34392_ (.A1(_10491_),
    .A2(_10496_),
    .ZN(_10540_));
 AOI21_X1 _34393_ (.A(_10540_),
    .B1(_10502_),
    .B2(_10521_),
    .ZN(_10541_));
 NOR2_X1 _34394_ (.A1(_10483_),
    .A2(_10464_),
    .ZN(_10542_));
 AOI211_X2 _34395_ (.A(_10539_),
    .B(_10541_),
    .C1(_10542_),
    .C2(_10482_),
    .ZN(_10543_));
 XNOR2_X2 _34396_ (.A(_10469_),
    .B(_10543_),
    .ZN(_10544_));
 OR2_X1 _34397_ (.A1(_10474_),
    .A2(_10464_),
    .ZN(_10545_));
 INV_X1 _34398_ (.A(_20459_),
    .ZN(_10546_));
 AOI21_X1 _34399_ (.A(_10545_),
    .B1(_10481_),
    .B2(_10546_),
    .ZN(_10547_));
 NOR2_X1 _34400_ (.A1(_20439_),
    .A2(_10491_),
    .ZN(_10548_));
 NOR2_X1 _34401_ (.A1(_10520_),
    .A2(_10519_),
    .ZN(_10549_));
 OAI21_X1 _34402_ (.A(_10474_),
    .B1(_20456_),
    .B2(_10549_),
    .ZN(_10550_));
 AOI221_X2 _34403_ (.A(_10547_),
    .B1(_10548_),
    .B2(_10550_),
    .C1(_20442_),
    .C2(_10492_),
    .ZN(_10551_));
 XOR2_X2 _34404_ (.A(_10473_),
    .B(_10551_),
    .Z(_10552_));
 AOI21_X1 _34405_ (.A(_20432_),
    .B1(_10502_),
    .B2(_10500_),
    .ZN(_10553_));
 MUX2_X2 _34406_ (.A(_10553_),
    .B(_10513_),
    .S(_10491_),
    .Z(_10554_));
 XNOR2_X2 _34407_ (.A(_20426_),
    .B(_10554_),
    .ZN(_10555_));
 AOI21_X2 _34408_ (.A(_10544_),
    .B1(_10552_),
    .B2(_10555_),
    .ZN(_10556_));
 MUX2_X2 _34409_ (.A(_10505_),
    .B(_10514_),
    .S(_10492_),
    .Z(_10557_));
 XNOR2_X2 _34410_ (.A(_20412_),
    .B(_10557_),
    .ZN(_10558_));
 OAI21_X2 _34411_ (.A(_10537_),
    .B1(_10556_),
    .B2(_10558_),
    .ZN(_10559_));
 NOR2_X1 _34412_ (.A1(_10527_),
    .A2(_10559_),
    .ZN(_10560_));
 NAND2_X2 _34413_ (.A1(_10457_),
    .A2(_10490_),
    .ZN(_10561_));
 OAI21_X2 _34414_ (.A(_10560_),
    .B1(_10561_),
    .B2(_10430_),
    .ZN(_10562_));
 OAI211_X2 _34415_ (.A(_10380_),
    .B(_10454_),
    .C1(_10425_),
    .C2(_10428_),
    .ZN(_10563_));
 NAND4_X4 _34416_ (.A1(_10365_),
    .A2(_10375_),
    .A3(_10411_),
    .A4(_10436_),
    .ZN(_10564_));
 NAND2_X1 _34417_ (.A1(_10382_),
    .A2(_10337_),
    .ZN(_10565_));
 OAI222_X2 _34418_ (.A1(_10384_),
    .A2(_10397_),
    .B1(_10398_),
    .B2(_10565_),
    .C1(_10432_),
    .C2(_10391_),
    .ZN(_10566_));
 OAI211_X4 _34419_ (.A(_10411_),
    .B(_10566_),
    .C1(_10425_),
    .C2(_10428_),
    .ZN(_10567_));
 XNOR2_X1 _34420_ (.A(_10486_),
    .B(_10557_),
    .ZN(_10568_));
 NOR2_X1 _34421_ (.A1(_20459_),
    .A2(_10464_),
    .ZN(_10569_));
 INV_X1 _34422_ (.A(_20456_),
    .ZN(_10570_));
 OAI21_X1 _34423_ (.A(_10570_),
    .B1(_10499_),
    .B2(_10477_),
    .ZN(_10571_));
 AOI22_X2 _34424_ (.A1(_10512_),
    .A2(_10569_),
    .B1(_10571_),
    .B2(_10464_),
    .ZN(_10572_));
 XNOR2_X2 _34425_ (.A(_10474_),
    .B(_10572_),
    .ZN(_10573_));
 INV_X2 _34426_ (.A(_10573_),
    .ZN(_10574_));
 NAND3_X4 _34427_ (.A1(_10568_),
    .A2(_10555_),
    .A3(_10574_),
    .ZN(_10575_));
 XOR2_X1 _34428_ (.A(_14494_),
    .B(_10498_),
    .Z(_10576_));
 XOR2_X1 _34429_ (.A(_14498_),
    .B(_10480_),
    .Z(_10577_));
 MUX2_X1 _34430_ (.A(_10576_),
    .B(_10577_),
    .S(_10492_),
    .Z(_10578_));
 CLKBUF_X3 _34431_ (.A(_10578_),
    .Z(_10579_));
 MUX2_X2 _34432_ (.A(_20463_),
    .B(_20465_),
    .S(_10492_),
    .Z(_10580_));
 NOR2_X1 _34433_ (.A1(_10579_),
    .A2(_10580_),
    .ZN(_10581_));
 NAND2_X1 _34434_ (.A1(_10492_),
    .A2(_10581_),
    .ZN(_10582_));
 NOR2_X1 _34435_ (.A1(_10575_),
    .A2(_10582_),
    .ZN(_10583_));
 NAND4_X1 _34436_ (.A1(_10563_),
    .A2(_10564_),
    .A3(_10567_),
    .A4(_10583_),
    .ZN(_10584_));
 INV_X1 _34437_ (.A(_10575_),
    .ZN(_10585_));
 NAND2_X1 _34438_ (.A1(_10465_),
    .A2(_10581_),
    .ZN(_10586_));
 AOI21_X2 _34439_ (.A(_10586_),
    .B1(_10331_),
    .B2(_10323_),
    .ZN(_10587_));
 NAND2_X1 _34440_ (.A1(_10585_),
    .A2(_10587_),
    .ZN(_10588_));
 AND2_X1 _34441_ (.A1(_10564_),
    .A2(_10567_),
    .ZN(_10589_));
 INV_X1 _34442_ (.A(_10498_),
    .ZN(_10590_));
 AOI21_X1 _34443_ (.A(_20401_),
    .B1(_14491_),
    .B2(_20402_),
    .ZN(_10591_));
 NOR2_X1 _34444_ (.A1(_10590_),
    .A2(_10591_),
    .ZN(_10592_));
 OAI21_X1 _34445_ (.A(_10464_),
    .B1(_10592_),
    .B2(_20407_),
    .ZN(_10593_));
 INV_X1 _34446_ (.A(_20452_),
    .ZN(_10594_));
 OAI21_X1 _34447_ (.A(_10480_),
    .B1(_10478_),
    .B2(_20403_),
    .ZN(_10595_));
 NAND2_X1 _34448_ (.A1(_10594_),
    .A2(_10595_),
    .ZN(_10596_));
 OAI21_X1 _34449_ (.A(_10593_),
    .B1(_10596_),
    .B2(_10464_),
    .ZN(_10597_));
 XNOR2_X2 _34450_ (.A(_10477_),
    .B(_10597_),
    .ZN(_10598_));
 MUX2_X2 _34451_ (.A(_14499_),
    .B(_14495_),
    .S(_10465_),
    .Z(_10599_));
 NOR2_X1 _34452_ (.A1(_10579_),
    .A2(_10599_),
    .ZN(_10600_));
 NOR2_X2 _34453_ (.A1(_10598_),
    .A2(_10600_),
    .ZN(_10601_));
 INV_X1 _34454_ (.A(_10601_),
    .ZN(_10602_));
 NOR3_X1 _34455_ (.A1(_20465_),
    .A2(_10465_),
    .A3(_10579_),
    .ZN(_10603_));
 NOR2_X1 _34456_ (.A1(_10419_),
    .A2(_10420_),
    .ZN(_10604_));
 NAND3_X1 _34457_ (.A1(_10377_),
    .A2(_10378_),
    .A3(_10454_),
    .ZN(_10605_));
 AOI21_X1 _34458_ (.A(_10605_),
    .B1(_10375_),
    .B2(_10365_),
    .ZN(_10606_));
 AOI221_X2 _34459_ (.A(_10602_),
    .B1(_10603_),
    .B2(_10604_),
    .C1(_10587_),
    .C2(_10606_),
    .ZN(_10607_));
 OAI221_X2 _34460_ (.A(_10584_),
    .B1(_10588_),
    .B2(_10589_),
    .C1(_10607_),
    .C2(_10575_),
    .ZN(_10608_));
 BUF_X4 _34461_ (.A(_10608_),
    .Z(_10609_));
 NOR2_X1 _34462_ (.A1(_10562_),
    .A2(_10609_),
    .ZN(_10610_));
 NOR2_X1 _34463_ (.A1(_10531_),
    .A2(_10610_),
    .ZN(_20467_));
 INV_X1 _34464_ (.A(_20467_),
    .ZN(_20469_));
 INV_X2 _34465_ (.A(_20472_),
    .ZN(_10611_));
 NOR2_X2 _34466_ (.A1(_10527_),
    .A2(_10516_),
    .ZN(_10612_));
 NOR4_X4 _34467_ (.A1(_10573_),
    .A2(_10579_),
    .A3(_10598_),
    .A4(_10552_),
    .ZN(_10613_));
 INV_X1 _34468_ (.A(_10488_),
    .ZN(_10614_));
 XNOR2_X2 _34469_ (.A(_10614_),
    .B(_10536_),
    .ZN(_10615_));
 XNOR2_X2 _34470_ (.A(_10483_),
    .B(_10554_),
    .ZN(_10616_));
 OR2_X1 _34471_ (.A1(_10616_),
    .A2(_10544_),
    .ZN(_10617_));
 OR3_X1 _34472_ (.A1(_10558_),
    .A2(_10615_),
    .A3(_10617_),
    .ZN(_10618_));
 OAI221_X2 _34473_ (.A(_10612_),
    .B1(_10613_),
    .B2(_10618_),
    .C1(_10463_),
    .C2(_10429_),
    .ZN(_10619_));
 OR2_X1 _34474_ (.A1(_10490_),
    .A2(_10528_),
    .ZN(_10620_));
 NOR2_X1 _34475_ (.A1(_10613_),
    .A2(_10618_),
    .ZN(_10621_));
 OR4_X1 _34476_ (.A1(_10429_),
    .A2(_10463_),
    .A3(_10620_),
    .A4(_10621_),
    .ZN(_10622_));
 AND3_X1 _34477_ (.A1(_10611_),
    .A2(_10619_),
    .A3(_10622_),
    .ZN(_10623_));
 AOI21_X1 _34478_ (.A(_10611_),
    .B1(_10619_),
    .B2(_10622_),
    .ZN(_10624_));
 OR2_X1 _34479_ (.A1(_10623_),
    .A2(_10624_),
    .ZN(_10625_));
 BUF_X4 _34480_ (.A(_10625_),
    .Z(_10626_));
 INV_X4 _34481_ (.A(_10626_),
    .ZN(_20493_));
 OR3_X2 _34482_ (.A1(_10429_),
    .A2(_10463_),
    .A3(_10620_),
    .ZN(_10627_));
 OAI21_X2 _34483_ (.A(_10612_),
    .B1(_10463_),
    .B2(_10430_),
    .ZN(_10628_));
 AND2_X2 _34484_ (.A1(_10627_),
    .A2(_10628_),
    .ZN(_10629_));
 AND4_X1 _34485_ (.A1(_10365_),
    .A2(_10375_),
    .A3(_10411_),
    .A4(_10436_),
    .ZN(_10630_));
 MUX2_X1 _34486_ (.A(_10454_),
    .B(_10566_),
    .S(_10411_),
    .Z(_10631_));
 AOI221_X2 _34487_ (.A(_10492_),
    .B1(_10630_),
    .B2(_10332_),
    .C1(_10631_),
    .C2(_10437_),
    .ZN(_10632_));
 NAND3_X1 _34488_ (.A1(_10257_),
    .A2(_10267_),
    .A3(_10453_),
    .ZN(_10633_));
 OAI21_X1 _34489_ (.A(_10633_),
    .B1(_10449_),
    .B2(_10273_),
    .ZN(_10634_));
 NAND3_X1 _34490_ (.A1(_10377_),
    .A2(_10378_),
    .A3(_10634_),
    .ZN(_10635_));
 OAI221_X2 _34491_ (.A(_10635_),
    .B1(_10566_),
    .B2(_10380_),
    .C1(_10425_),
    .C2(_10428_),
    .ZN(_10636_));
 AOI211_X2 _34492_ (.A(_10604_),
    .B(_10465_),
    .C1(_10564_),
    .C2(_10636_),
    .ZN(_10637_));
 NOR2_X2 _34493_ (.A1(_10632_),
    .A2(_10637_),
    .ZN(_10638_));
 BUF_X4 _34494_ (.A(_20468_),
    .Z(_10639_));
 OAI21_X1 _34495_ (.A(_10629_),
    .B1(_10638_),
    .B2(_10639_),
    .ZN(_10640_));
 AOI21_X4 _34496_ (.A(_10528_),
    .B1(_10457_),
    .B2(_10437_),
    .ZN(_10641_));
 NOR2_X2 _34497_ (.A1(_10558_),
    .A2(_10556_),
    .ZN(_10642_));
 NOR2_X4 _34498_ (.A1(_10642_),
    .A2(_10615_),
    .ZN(_10643_));
 NOR3_X4 _34499_ (.A1(_10429_),
    .A2(_10463_),
    .A3(_10516_),
    .ZN(_10644_));
 BUF_X1 _34500_ (.A(_14506_),
    .Z(_10645_));
 INV_X2 _34501_ (.A(_10645_),
    .ZN(_14501_));
 NOR2_X1 _34502_ (.A1(_14501_),
    .A2(_10527_),
    .ZN(_10646_));
 OAI21_X4 _34503_ (.A(_10646_),
    .B1(_10561_),
    .B2(_10429_),
    .ZN(_10647_));
 NOR4_X2 _34504_ (.A1(_10641_),
    .A2(_10643_),
    .A3(_10644_),
    .A4(_10647_),
    .ZN(_10648_));
 NOR3_X2 _34505_ (.A1(_10647_),
    .A2(_10632_),
    .A3(_10637_),
    .ZN(_10649_));
 NOR3_X1 _34506_ (.A1(_10641_),
    .A2(_10644_),
    .A3(_10647_),
    .ZN(_10650_));
 AOI211_X2 _34507_ (.A(_10648_),
    .B(_10649_),
    .C1(_10609_),
    .C2(_10650_),
    .ZN(_10651_));
 NOR3_X1 _34508_ (.A1(_20463_),
    .A2(_10492_),
    .A3(_10579_),
    .ZN(_10652_));
 OAI21_X2 _34509_ (.A(_10652_),
    .B1(_10420_),
    .B2(net343),
    .ZN(_10653_));
 OAI221_X2 _34510_ (.A(_10601_),
    .B1(_10582_),
    .B2(_10332_),
    .C1(_10653_),
    .C2(_10563_),
    .ZN(_10654_));
 AOI21_X2 _34511_ (.A(_10653_),
    .B1(_10564_),
    .B2(_10567_),
    .ZN(_10655_));
 AND3_X1 _34512_ (.A1(_10603_),
    .A2(_10564_),
    .A3(_10636_),
    .ZN(_10656_));
 NAND2_X1 _34513_ (.A1(_10568_),
    .A2(_10537_),
    .ZN(_10657_));
 NOR2_X2 _34514_ (.A1(_10617_),
    .A2(_10657_),
    .ZN(_10658_));
 XNOR2_X2 _34515_ (.A(_10473_),
    .B(_10551_),
    .ZN(_10659_));
 NAND2_X1 _34516_ (.A1(_10574_),
    .A2(_10659_),
    .ZN(_10660_));
 AND2_X1 _34517_ (.A1(_20463_),
    .A2(_10465_),
    .ZN(_10661_));
 AOI21_X2 _34518_ (.A(_10661_),
    .B1(_10492_),
    .B2(_20465_),
    .ZN(_10662_));
 NAND2_X1 _34519_ (.A1(_10662_),
    .A2(_10599_),
    .ZN(_10663_));
 NOR2_X1 _34520_ (.A1(_10579_),
    .A2(_10598_),
    .ZN(_10664_));
 AOI21_X1 _34521_ (.A(_10660_),
    .B1(_10663_),
    .B2(_10664_),
    .ZN(_10665_));
 NAND2_X1 _34522_ (.A1(_10658_),
    .A2(_10665_),
    .ZN(_10666_));
 OR4_X1 _34523_ (.A1(_10654_),
    .A2(_10655_),
    .A3(_10656_),
    .A4(_10666_),
    .ZN(_10667_));
 NOR2_X1 _34524_ (.A1(_10611_),
    .A2(_10621_),
    .ZN(_10668_));
 AOI221_X2 _34525_ (.A(_10668_),
    .B1(_10628_),
    .B2(_10627_),
    .C1(_10611_),
    .C2(_10658_),
    .ZN(_10669_));
 NAND2_X1 _34526_ (.A1(_10667_),
    .A2(_10669_),
    .ZN(_10670_));
 OAI21_X1 _34527_ (.A(_10640_),
    .B1(_10651_),
    .B2(_10670_),
    .ZN(_10671_));
 BUF_X4 _34528_ (.A(_10629_),
    .Z(_10672_));
 NAND3_X1 _34529_ (.A1(_10639_),
    .A2(_10672_),
    .A3(_10662_),
    .ZN(_10673_));
 NAND2_X1 _34530_ (.A1(_10671_),
    .A2(_10673_),
    .ZN(_10674_));
 INV_X4 _34531_ (.A(_20468_),
    .ZN(_10675_));
 NAND2_X1 _34532_ (.A1(_10675_),
    .A2(_10580_),
    .ZN(_10676_));
 OAI21_X2 _34533_ (.A(_10676_),
    .B1(_10599_),
    .B2(_10675_),
    .ZN(_10677_));
 OAI211_X2 _34534_ (.A(_10650_),
    .B(_10638_),
    .C1(_10642_),
    .C2(_10609_),
    .ZN(_10678_));
 NOR2_X1 _34535_ (.A1(_14501_),
    .A2(_10580_),
    .ZN(_10679_));
 NAND2_X1 _34536_ (.A1(_10465_),
    .A2(_10526_),
    .ZN(_10680_));
 OAI21_X2 _34537_ (.A(_10680_),
    .B1(_10561_),
    .B2(_10430_),
    .ZN(_10681_));
 NOR2_X1 _34538_ (.A1(_10681_),
    .A2(_10559_),
    .ZN(_10682_));
 AND4_X1 _34539_ (.A1(_10563_),
    .A2(_10564_),
    .A3(_10567_),
    .A4(_10583_),
    .ZN(_10683_));
 NOR2_X1 _34540_ (.A1(_10575_),
    .A2(_10653_),
    .ZN(_10684_));
 NAND2_X1 _34541_ (.A1(_10564_),
    .A2(_10567_),
    .ZN(_10685_));
 AOI221_X4 _34542_ (.A(_10683_),
    .B1(_10684_),
    .B2(_10685_),
    .C1(_10654_),
    .C2(_10585_),
    .ZN(_10686_));
 NAND2_X1 _34543_ (.A1(_10682_),
    .A2(_10686_),
    .ZN(_10687_));
 OAI21_X4 _34544_ (.A(_10516_),
    .B1(_10463_),
    .B2(_10429_),
    .ZN(_10688_));
 NAND3_X4 _34545_ (.A1(_10437_),
    .A2(_10457_),
    .A3(_10528_),
    .ZN(_10689_));
 NAND2_X4 _34546_ (.A1(_10688_),
    .A2(_10689_),
    .ZN(_10690_));
 NAND2_X1 _34547_ (.A1(_10645_),
    .A2(_10662_),
    .ZN(_10691_));
 NOR4_X1 _34548_ (.A1(_14501_),
    .A2(_10641_),
    .A3(_10537_),
    .A4(_10644_),
    .ZN(_10692_));
 AOI22_X1 _34549_ (.A1(_10690_),
    .A2(_10691_),
    .B1(_10692_),
    .B2(_10638_),
    .ZN(_10693_));
 BUF_X4 _34550_ (.A(_10681_),
    .Z(_10694_));
 OAI221_X2 _34551_ (.A(_10678_),
    .B1(_10679_),
    .B2(_10687_),
    .C1(_10693_),
    .C2(_10694_),
    .ZN(_10695_));
 AND2_X2 _34552_ (.A1(_10667_),
    .A2(_10669_),
    .ZN(_10696_));
 AOI22_X4 _34553_ (.A1(_10672_),
    .A2(_10677_),
    .B1(_10695_),
    .B2(_10696_),
    .ZN(_10697_));
 NOR2_X1 _34554_ (.A1(_10674_),
    .A2(_10697_),
    .ZN(_20474_));
 NOR2_X4 _34555_ (.A1(net344),
    .A2(_10231_),
    .ZN(_10698_));
 AOI22_X4 _34556_ (.A1(\g_reduce0[0].adder.b[0] ),
    .A2(net344),
    .B1(_10698_),
    .B2(\g_reduce0[0].adder.a[0] ),
    .ZN(_10699_));
 OR4_X4 _34557_ (.A1(\g_reduce0[0].adder.a[11] ),
    .A2(_10224_),
    .A3(_10225_),
    .A4(_10226_),
    .ZN(_10700_));
 NAND2_X2 _34558_ (.A1(_10700_),
    .A2(_10231_),
    .ZN(_10701_));
 INV_X1 _34559_ (.A(_20477_),
    .ZN(_10702_));
 NAND2_X4 _34560_ (.A1(_10627_),
    .A2(_10628_),
    .ZN(_10703_));
 NOR4_X4 _34561_ (.A1(_10654_),
    .A2(_10655_),
    .A3(_10656_),
    .A4(_10666_),
    .ZN(_10704_));
 AND2_X1 _34562_ (.A1(_10613_),
    .A2(_10658_),
    .ZN(_10705_));
 OR2_X1 _34563_ (.A1(_10681_),
    .A2(_10705_),
    .ZN(_10706_));
 OAI22_X4 _34564_ (.A1(_10694_),
    .A2(_10703_),
    .B1(_10704_),
    .B2(_10706_),
    .ZN(_20497_));
 AND3_X1 _34565_ (.A1(_20470_),
    .A2(_20493_),
    .A3(_20497_),
    .ZN(_10707_));
 OAI21_X1 _34566_ (.A(_10697_),
    .B1(_10707_),
    .B2(_10672_),
    .ZN(_10708_));
 MUX2_X1 _34567_ (.A(_10708_),
    .B(_10697_),
    .S(_10674_),
    .Z(_10709_));
 NOR3_X4 _34568_ (.A1(_10629_),
    .A2(_10704_),
    .A3(_10705_),
    .ZN(_10710_));
 NOR3_X2 _34569_ (.A1(_10641_),
    .A2(_10537_),
    .A3(_10644_),
    .ZN(_10711_));
 AOI21_X1 _34570_ (.A(_10616_),
    .B1(_10537_),
    .B2(_10558_),
    .ZN(_10712_));
 INV_X1 _34571_ (.A(_10712_),
    .ZN(_10713_));
 OAI22_X4 _34572_ (.A1(_10544_),
    .A2(_10711_),
    .B1(_10713_),
    .B2(_10690_),
    .ZN(_10714_));
 OR3_X1 _34573_ (.A1(_20493_),
    .A2(_10647_),
    .A3(_10714_),
    .ZN(_10715_));
 NOR2_X1 _34574_ (.A1(_10694_),
    .A2(_10537_),
    .ZN(_10716_));
 OAI21_X1 _34575_ (.A(_10716_),
    .B1(_10690_),
    .B2(_10558_),
    .ZN(_10717_));
 NOR3_X2 _34576_ (.A1(_10641_),
    .A2(_10643_),
    .A3(_10644_),
    .ZN(_10718_));
 NAND2_X1 _34577_ (.A1(_10575_),
    .A2(_10643_),
    .ZN(_10719_));
 NAND3_X2 _34578_ (.A1(_10688_),
    .A2(_10689_),
    .A3(_10719_),
    .ZN(_10720_));
 AOI22_X4 _34579_ (.A1(_10573_),
    .A2(_10718_),
    .B1(_10720_),
    .B2(_10552_),
    .ZN(_10721_));
 MUX2_X1 _34580_ (.A(_10717_),
    .B(_10721_),
    .S(_10626_),
    .Z(_10722_));
 CLKBUF_X3 _34581_ (.A(_10645_),
    .Z(_10723_));
 OAI21_X1 _34582_ (.A(_10715_),
    .B1(_10722_),
    .B2(_10723_),
    .ZN(_10724_));
 NOR2_X1 _34583_ (.A1(_20497_),
    .A2(_10690_),
    .ZN(_10725_));
 AND2_X1 _34584_ (.A1(_10609_),
    .A2(_10650_),
    .ZN(_10726_));
 OR3_X2 _34585_ (.A1(_10726_),
    .A2(_10648_),
    .A3(_10649_),
    .ZN(_10727_));
 INV_X1 _34586_ (.A(_10579_),
    .ZN(_10728_));
 NAND2_X1 _34587_ (.A1(_10645_),
    .A2(_10728_),
    .ZN(_10729_));
 NAND2_X1 _34588_ (.A1(_14501_),
    .A2(_10662_),
    .ZN(_10730_));
 AOI221_X2 _34589_ (.A(_10690_),
    .B1(_10729_),
    .B2(_10730_),
    .C1(_10686_),
    .C2(_10643_),
    .ZN(_10731_));
 NOR2_X4 _34590_ (.A1(_10641_),
    .A2(_10644_),
    .ZN(_10732_));
 OAI21_X4 _34591_ (.A(_10732_),
    .B1(_10609_),
    .B2(_10559_),
    .ZN(_10733_));
 NAND2_X1 _34592_ (.A1(_10645_),
    .A2(_10598_),
    .ZN(_10734_));
 OAI21_X1 _34593_ (.A(_10734_),
    .B1(_10599_),
    .B2(_10645_),
    .ZN(_10735_));
 INV_X1 _34594_ (.A(_10735_),
    .ZN(_10736_));
 AOI211_X2 _34595_ (.A(_10694_),
    .B(_10731_),
    .C1(_10733_),
    .C2(_10736_),
    .ZN(_10737_));
 MUX2_X1 _34596_ (.A(_10727_),
    .B(_10737_),
    .S(_20493_),
    .Z(_10738_));
 AOI221_X2 _34597_ (.A(_10694_),
    .B1(_10710_),
    .B2(_10724_),
    .C1(_10725_),
    .C2(_10738_),
    .ZN(_10739_));
 AOI21_X4 _34598_ (.A(_10739_),
    .B1(_10672_),
    .B2(_10639_),
    .ZN(_10740_));
 MUX2_X1 _34599_ (.A(_10694_),
    .B(_10690_),
    .S(_10675_),
    .Z(_10741_));
 NOR3_X1 _34600_ (.A1(_10672_),
    .A2(_20493_),
    .A3(_20497_),
    .ZN(_10742_));
 AND2_X1 _34601_ (.A1(_10626_),
    .A2(_10710_),
    .ZN(_10743_));
 MUX2_X1 _34602_ (.A(_10555_),
    .B(_10574_),
    .S(_14501_),
    .Z(_10744_));
 INV_X1 _34603_ (.A(_10744_),
    .ZN(_10745_));
 NOR2_X1 _34604_ (.A1(_10562_),
    .A2(_10745_),
    .ZN(_10746_));
 NOR4_X2 _34605_ (.A1(_10430_),
    .A2(_10463_),
    .A3(_10490_),
    .A4(_10516_),
    .ZN(_10747_));
 AOI221_X2 _34606_ (.A(_10528_),
    .B1(_10526_),
    .B2(_10465_),
    .C1(_10437_),
    .C2(_10457_),
    .ZN(_10748_));
 NOR2_X1 _34607_ (.A1(_10645_),
    .A2(_10598_),
    .ZN(_10749_));
 AOI21_X1 _34608_ (.A(_10749_),
    .B1(_10659_),
    .B2(_10645_),
    .ZN(_10750_));
 NOR3_X1 _34609_ (.A1(_10747_),
    .A2(_10748_),
    .A3(_10750_),
    .ZN(_10751_));
 MUX2_X1 _34610_ (.A(_10746_),
    .B(_10751_),
    .S(_10609_),
    .Z(_10752_));
 OAI21_X1 _34611_ (.A(_10744_),
    .B1(_10748_),
    .B2(_10747_),
    .ZN(_10753_));
 INV_X1 _34612_ (.A(_10750_),
    .ZN(_10754_));
 NAND2_X1 _34613_ (.A1(_10562_),
    .A2(_10754_),
    .ZN(_10755_));
 OAI21_X1 _34614_ (.A(_10753_),
    .B1(_10755_),
    .B2(_10531_),
    .ZN(_10756_));
 NOR2_X1 _34615_ (.A1(_10752_),
    .A2(_10756_),
    .ZN(_10757_));
 AOI221_X1 _34616_ (.A(_10741_),
    .B1(_10742_),
    .B2(_20470_),
    .C1(_10743_),
    .C2(_10757_),
    .ZN(_10758_));
 OR3_X1 _34617_ (.A1(_10728_),
    .A2(_10562_),
    .A3(_10647_),
    .ZN(_10759_));
 OR4_X1 _34618_ (.A1(_10641_),
    .A2(_10599_),
    .A3(_10644_),
    .A4(_10647_),
    .ZN(_10760_));
 MUX2_X1 _34619_ (.A(_10759_),
    .B(_10760_),
    .S(_10609_),
    .Z(_10761_));
 NOR2_X1 _34620_ (.A1(_14501_),
    .A2(_10681_),
    .ZN(_10762_));
 AOI21_X2 _34621_ (.A(_10728_),
    .B1(_10530_),
    .B2(_10517_),
    .ZN(_10763_));
 NOR4_X2 _34622_ (.A1(_10641_),
    .A2(_10599_),
    .A3(_10643_),
    .A4(_10644_),
    .ZN(_10764_));
 OAI21_X2 _34623_ (.A(_10762_),
    .B1(_10763_),
    .B2(_10764_),
    .ZN(_10765_));
 OR2_X1 _34624_ (.A1(_10580_),
    .A2(_10562_),
    .ZN(_10766_));
 OAI22_X4 _34625_ (.A1(_10580_),
    .A2(_10732_),
    .B1(_10766_),
    .B2(_10609_),
    .ZN(_10767_));
 NOR2_X1 _34626_ (.A1(_10723_),
    .A2(_10694_),
    .ZN(_10768_));
 OAI21_X1 _34627_ (.A(_10643_),
    .B1(_10601_),
    .B2(_10575_),
    .ZN(_10769_));
 NAND3_X1 _34628_ (.A1(_10688_),
    .A2(_10689_),
    .A3(_10769_),
    .ZN(_10770_));
 OAI21_X2 _34629_ (.A(_10768_),
    .B1(_10770_),
    .B2(_10638_),
    .ZN(_10771_));
 OAI211_X4 _34630_ (.A(_10761_),
    .B(_10765_),
    .C1(_10767_),
    .C2(_10771_),
    .ZN(_10772_));
 NOR3_X2 _34631_ (.A1(_10672_),
    .A2(_10626_),
    .A3(_20497_),
    .ZN(_10773_));
 NAND3_X1 _34632_ (.A1(_10688_),
    .A2(_10544_),
    .A3(_10689_),
    .ZN(_10774_));
 OAI21_X1 _34633_ (.A(_10774_),
    .B1(_10711_),
    .B2(_10568_),
    .ZN(_10775_));
 NAND2_X1 _34634_ (.A1(_10537_),
    .A2(_10732_),
    .ZN(_10776_));
 MUX2_X1 _34635_ (.A(_10775_),
    .B(_10776_),
    .S(_10723_),
    .Z(_10777_));
 NOR2_X1 _34636_ (.A1(_10672_),
    .A2(_10626_),
    .ZN(_10778_));
 AOI22_X1 _34637_ (.A1(_10772_),
    .A2(_10773_),
    .B1(_10777_),
    .B2(_10778_),
    .ZN(_10779_));
 AND2_X1 _34638_ (.A1(_10758_),
    .A2(_10779_),
    .ZN(_10780_));
 NAND3_X1 _34639_ (.A1(_10688_),
    .A2(_10689_),
    .A3(_10679_),
    .ZN(_10781_));
 AOI21_X1 _34640_ (.A(_10781_),
    .B1(_10686_),
    .B2(_10643_),
    .ZN(_10782_));
 NAND2_X1 _34641_ (.A1(_10723_),
    .A2(_10599_),
    .ZN(_10783_));
 OAI21_X1 _34642_ (.A(_10783_),
    .B1(_10638_),
    .B2(_10723_),
    .ZN(_10784_));
 AOI21_X2 _34643_ (.A(_10782_),
    .B1(_10784_),
    .B2(_10733_),
    .ZN(_10785_));
 AND2_X1 _34644_ (.A1(_10785_),
    .A2(_10773_),
    .ZN(_10786_));
 NAND2_X1 _34645_ (.A1(_10733_),
    .A2(_10749_),
    .ZN(_10787_));
 NAND2_X1 _34646_ (.A1(_10723_),
    .A2(_10721_),
    .ZN(_10788_));
 OR3_X1 _34647_ (.A1(_10723_),
    .A2(_10579_),
    .A3(_10733_),
    .ZN(_10789_));
 AND4_X1 _34648_ (.A1(_10743_),
    .A2(_10787_),
    .A3(_10788_),
    .A4(_10789_),
    .ZN(_10790_));
 NOR2_X1 _34649_ (.A1(_14501_),
    .A2(_10717_),
    .ZN(_10791_));
 NOR2_X1 _34650_ (.A1(_10723_),
    .A2(_10714_),
    .ZN(_10792_));
 OAI21_X1 _34651_ (.A(_10778_),
    .B1(_10791_),
    .B2(_10792_),
    .ZN(_10793_));
 MUX2_X1 _34652_ (.A(_10537_),
    .B(_10732_),
    .S(_10639_),
    .Z(_10794_));
 CLKBUF_X3 _34653_ (.A(_10703_),
    .Z(_10795_));
 OAI21_X2 _34654_ (.A(_10793_),
    .B1(_10794_),
    .B2(_10795_),
    .ZN(_10796_));
 NOR3_X2 _34655_ (.A1(_10786_),
    .A2(_10790_),
    .A3(_10796_),
    .ZN(_10797_));
 NOR2_X1 _34656_ (.A1(_10780_),
    .A2(_10797_),
    .ZN(_10798_));
 INV_X1 _34657_ (.A(_20470_),
    .ZN(_10799_));
 OAI33_X1 _34658_ (.A1(_10799_),
    .A2(_10623_),
    .A3(_10624_),
    .B1(_10704_),
    .B2(_10705_),
    .B3(_10694_),
    .ZN(_10800_));
 MUX2_X1 _34659_ (.A(_10616_),
    .B(_10544_),
    .S(_10639_),
    .Z(_10801_));
 MUX2_X1 _34660_ (.A(_10800_),
    .B(_10801_),
    .S(_10629_),
    .Z(_10802_));
 NAND2_X1 _34661_ (.A1(_10626_),
    .A2(_10710_),
    .ZN(_10803_));
 NOR3_X1 _34662_ (.A1(_10694_),
    .A2(_10752_),
    .A3(_10756_),
    .ZN(_10804_));
 OAI221_X2 _34663_ (.A(_10802_),
    .B1(_10772_),
    .B2(_10803_),
    .C1(_10670_),
    .C2(_10804_),
    .ZN(_10805_));
 MUX2_X1 _34664_ (.A(_10558_),
    .B(_10544_),
    .S(_10675_),
    .Z(_10806_));
 AOI22_X2 _34665_ (.A1(_10672_),
    .A2(_10806_),
    .B1(_10773_),
    .B2(_10727_),
    .ZN(_10807_));
 OAI221_X2 _34666_ (.A(_20493_),
    .B1(_10647_),
    .B2(_10714_),
    .C1(_10721_),
    .C2(_10723_),
    .ZN(_10808_));
 OAI211_X2 _34667_ (.A(_10710_),
    .B(_10808_),
    .C1(_10737_),
    .C2(_20493_),
    .ZN(_10809_));
 AOI21_X1 _34668_ (.A(_10805_),
    .B1(_10807_),
    .B2(_10809_),
    .ZN(_10810_));
 XNOR2_X1 _34669_ (.A(_20472_),
    .B(_10664_),
    .ZN(_10811_));
 NOR2_X1 _34670_ (.A1(_10430_),
    .A2(_10561_),
    .ZN(_10812_));
 NOR2_X1 _34671_ (.A1(_10527_),
    .A2(_10812_),
    .ZN(_10813_));
 AOI221_X1 _34672_ (.A(_10611_),
    .B1(_10813_),
    .B2(_10629_),
    .C1(_10682_),
    .C2(_10686_),
    .ZN(_10814_));
 NOR3_X1 _34673_ (.A1(_10660_),
    .A2(_10811_),
    .A3(_10814_),
    .ZN(_10815_));
 NAND4_X1 _34674_ (.A1(_10703_),
    .A2(_10658_),
    .A3(_10695_),
    .A4(_10815_),
    .ZN(_10816_));
 OR2_X1 _34675_ (.A1(_10645_),
    .A2(_10681_),
    .ZN(_10817_));
 NOR3_X1 _34676_ (.A1(_10641_),
    .A2(_10552_),
    .A3(_10644_),
    .ZN(_10818_));
 OR3_X1 _34677_ (.A1(_10645_),
    .A2(_10681_),
    .A3(_10559_),
    .ZN(_10819_));
 OAI22_X1 _34678_ (.A1(_10817_),
    .A2(_10818_),
    .B1(_10819_),
    .B2(_10609_),
    .ZN(_10820_));
 NOR2_X1 _34679_ (.A1(_10616_),
    .A2(_10562_),
    .ZN(_10821_));
 AOI22_X1 _34680_ (.A1(_10531_),
    .A2(_10555_),
    .B1(_10686_),
    .B2(_10821_),
    .ZN(_10822_));
 AOI221_X1 _34681_ (.A(_10626_),
    .B1(_10762_),
    .B2(_10775_),
    .C1(_10820_),
    .C2(_10822_),
    .ZN(_10823_));
 OR4_X1 _34682_ (.A1(_10672_),
    .A2(_10704_),
    .A3(_10705_),
    .A4(_10823_),
    .ZN(_10824_));
 OR4_X1 _34683_ (.A1(_14501_),
    .A2(_10694_),
    .A3(_10574_),
    .A4(_10718_),
    .ZN(_10825_));
 NAND4_X1 _34684_ (.A1(_10723_),
    .A2(_10813_),
    .A3(_10703_),
    .A4(_10598_),
    .ZN(_10826_));
 OAI21_X1 _34685_ (.A(_10825_),
    .B1(_10826_),
    .B2(_10610_),
    .ZN(_10827_));
 NOR2_X1 _34686_ (.A1(_10763_),
    .A2(_10764_),
    .ZN(_10828_));
 OR3_X1 _34687_ (.A1(_10641_),
    .A2(_10599_),
    .A3(_10644_),
    .ZN(_10829_));
 OR2_X1 _34688_ (.A1(_10728_),
    .A2(_10562_),
    .ZN(_10830_));
 MUX2_X1 _34689_ (.A(_10829_),
    .B(_10830_),
    .S(_10686_),
    .Z(_10831_));
 AOI21_X2 _34690_ (.A(_10817_),
    .B1(_10828_),
    .B2(_10831_),
    .ZN(_10832_));
 NOR3_X1 _34691_ (.A1(_20493_),
    .A2(_10827_),
    .A3(_10832_),
    .ZN(_10833_));
 MUX2_X1 _34692_ (.A(_10568_),
    .B(_10537_),
    .S(_10639_),
    .Z(_10834_));
 OAI221_X2 _34693_ (.A(_10816_),
    .B1(_10824_),
    .B2(_10833_),
    .C1(_10834_),
    .C2(_10703_),
    .ZN(_10835_));
 NAND2_X1 _34694_ (.A1(_10810_),
    .A2(_10835_),
    .ZN(_10836_));
 XNOR2_X1 _34695_ (.A(_10611_),
    .B(_10621_),
    .ZN(_10837_));
 AND3_X1 _34696_ (.A1(_20470_),
    .A2(_10710_),
    .A3(_10837_),
    .ZN(_10838_));
 MUX2_X1 _34697_ (.A(_10579_),
    .B(_10598_),
    .S(_10639_),
    .Z(_10839_));
 AOI221_X2 _34698_ (.A(_10838_),
    .B1(_10839_),
    .B2(_10672_),
    .C1(_10772_),
    .C2(_10696_),
    .ZN(_10840_));
 INV_X1 _34699_ (.A(_10840_),
    .ZN(_10841_));
 MUX2_X1 _34700_ (.A(_10573_),
    .B(_10598_),
    .S(_10675_),
    .Z(_10842_));
 AOI222_X2 _34701_ (.A1(_10696_),
    .A2(_10737_),
    .B1(_10743_),
    .B2(_10727_),
    .C1(_10842_),
    .C2(_10629_),
    .ZN(_10843_));
 MUX2_X1 _34702_ (.A(_10728_),
    .B(_10599_),
    .S(_10675_),
    .Z(_10844_));
 NOR2_X1 _34703_ (.A1(_10703_),
    .A2(_10844_),
    .ZN(_10845_));
 AOI21_X2 _34704_ (.A(_10845_),
    .B1(_10785_),
    .B2(_10696_),
    .ZN(_10846_));
 NOR4_X2 _34705_ (.A1(_10674_),
    .A2(_10697_),
    .A3(_10843_),
    .A4(_10846_),
    .ZN(_10847_));
 MUX2_X1 _34706_ (.A(_10574_),
    .B(_10659_),
    .S(_10639_),
    .Z(_10848_));
 NOR3_X2 _34707_ (.A1(_10626_),
    .A2(_10827_),
    .A3(_10832_),
    .ZN(_10849_));
 OAI21_X2 _34708_ (.A(_10710_),
    .B1(_10695_),
    .B2(_20493_),
    .ZN(_10850_));
 OAI22_X4 _34709_ (.A1(_10703_),
    .A2(_10848_),
    .B1(_10849_),
    .B2(_10850_),
    .ZN(_10851_));
 MUX2_X1 _34710_ (.A(_10679_),
    .B(_10784_),
    .S(_10733_),
    .Z(_10852_));
 NAND2_X1 _34711_ (.A1(_10696_),
    .A2(_10789_),
    .ZN(_10853_));
 NAND3_X1 _34712_ (.A1(_10813_),
    .A2(_10787_),
    .A3(_10788_),
    .ZN(_10854_));
 MUX2_X1 _34713_ (.A(_10555_),
    .B(_10659_),
    .S(_10675_),
    .Z(_10855_));
 OAI222_X2 _34714_ (.A1(_10803_),
    .A2(_10852_),
    .B1(_10853_),
    .B2(_10854_),
    .C1(_10855_),
    .C2(_10703_),
    .ZN(_10856_));
 NAND4_X1 _34715_ (.A1(_10841_),
    .A2(_10847_),
    .A3(_10851_),
    .A4(_10856_),
    .ZN(_10857_));
 NOR2_X1 _34716_ (.A1(_10836_),
    .A2(_10857_),
    .ZN(_10858_));
 AND2_X1 _34717_ (.A1(_10798_),
    .A2(_10858_),
    .ZN(_10859_));
 XNOR2_X2 _34718_ (.A(_10740_),
    .B(_10859_),
    .ZN(_10860_));
 MUX2_X1 _34719_ (.A(_10702_),
    .B(_10709_),
    .S(_10860_),
    .Z(_10861_));
 OAI21_X2 _34720_ (.A(_10699_),
    .B1(_10701_),
    .B2(_10861_),
    .ZN(_00000_));
 BUF_X4 _34721_ (.A(_10700_),
    .Z(_10862_));
 NOR4_X4 _34722_ (.A1(\g_reduce0[0].adder.b[11] ),
    .A2(\g_reduce0[0].adder.b[12] ),
    .A3(_10228_),
    .A4(_10229_),
    .ZN(_10863_));
 NAND2_X4 _34723_ (.A1(_10700_),
    .A2(_10863_),
    .ZN(_10864_));
 OAI22_X4 _34724_ (.A1(\g_reduce0[0].adder.b[1] ),
    .A2(_10862_),
    .B1(_10864_),
    .B2(\g_reduce0[0].adder.a[1] ),
    .ZN(_10865_));
 INV_X1 _34725_ (.A(_20476_),
    .ZN(_10866_));
 XNOR2_X1 _34726_ (.A(_10866_),
    .B(_10840_),
    .ZN(_10867_));
 MUX2_X1 _34727_ (.A(_10867_),
    .B(_10702_),
    .S(_10860_),
    .Z(_10868_));
 NOR2_X4 _34728_ (.A1(_10227_),
    .A2(_10863_),
    .ZN(_10869_));
 AOI21_X2 _34729_ (.A(_10865_),
    .B1(_10868_),
    .B2(_10869_),
    .ZN(_00007_));
 INV_X1 _34730_ (.A(_10846_),
    .ZN(_20475_));
 NAND3_X1 _34731_ (.A1(_20474_),
    .A2(_10841_),
    .A3(_20475_),
    .ZN(_10870_));
 XOR2_X1 _34732_ (.A(_10843_),
    .B(_10870_),
    .Z(_10871_));
 NAND2_X1 _34733_ (.A1(_10869_),
    .A2(_10871_),
    .ZN(_10872_));
 OR2_X1 _34734_ (.A1(_10701_),
    .A2(_10867_),
    .ZN(_10873_));
 MUX2_X1 _34735_ (.A(_10872_),
    .B(_10873_),
    .S(_10860_),
    .Z(_10874_));
 AOI22_X2 _34736_ (.A1(\g_reduce0[0].adder.b[2] ),
    .A2(net344),
    .B1(_10698_),
    .B2(\g_reduce0[0].adder.a[2] ),
    .ZN(_10875_));
 NAND2_X1 _34737_ (.A1(_10874_),
    .A2(_10875_),
    .ZN(_00008_));
 NOR3_X1 _34738_ (.A1(_10866_),
    .A2(_10843_),
    .A3(_10840_),
    .ZN(_10876_));
 XNOR2_X2 _34739_ (.A(_10851_),
    .B(_10876_),
    .ZN(_10877_));
 OR3_X1 _34740_ (.A1(_10860_),
    .A2(_10701_),
    .A3(_10877_),
    .ZN(_10878_));
 NOR2_X2 _34741_ (.A1(\g_reduce0[0].adder.b[3] ),
    .A2(_10862_),
    .ZN(_10879_));
 AOI21_X2 _34742_ (.A(net344),
    .B1(_10863_),
    .B2(\g_reduce0[0].adder.a[3] ),
    .ZN(_10880_));
 INV_X1 _34743_ (.A(_10860_),
    .ZN(_20480_));
 OAI221_X2 _34744_ (.A(_10878_),
    .B1(_10879_),
    .B2(_10880_),
    .C1(_10872_),
    .C2(_20480_),
    .ZN(_00009_));
 OAI22_X4 _34745_ (.A1(\g_reduce0[0].adder.b[4] ),
    .A2(_10862_),
    .B1(_10864_),
    .B2(\g_reduce0[0].adder.a[4] ),
    .ZN(_10881_));
 NOR3_X1 _34746_ (.A1(_10740_),
    .A2(_10859_),
    .A3(_10877_),
    .ZN(_10882_));
 INV_X2 _34747_ (.A(_10740_),
    .ZN(_10883_));
 AND3_X1 _34748_ (.A1(_10841_),
    .A2(_10847_),
    .A3(_10851_),
    .ZN(_10884_));
 NOR2_X1 _34749_ (.A1(_10856_),
    .A2(_10884_),
    .ZN(_10885_));
 NOR2_X1 _34750_ (.A1(_10883_),
    .A2(_10885_),
    .ZN(_10886_));
 AND2_X1 _34751_ (.A1(_10856_),
    .A2(_10884_),
    .ZN(_10887_));
 NAND2_X1 _34752_ (.A1(_10798_),
    .A2(_10858_),
    .ZN(_10888_));
 OAI21_X1 _34753_ (.A(_10887_),
    .B1(_10888_),
    .B2(_20476_),
    .ZN(_10889_));
 AOI21_X1 _34754_ (.A(_10882_),
    .B1(_10886_),
    .B2(_10889_),
    .ZN(_10890_));
 AOI21_X2 _34755_ (.A(_10881_),
    .B1(_10890_),
    .B2(_10869_),
    .ZN(_00010_));
 OAI22_X4 _34756_ (.A1(\g_reduce0[0].adder.b[5] ),
    .A2(_10862_),
    .B1(_10864_),
    .B2(\g_reduce0[0].adder.a[5] ),
    .ZN(_10891_));
 NAND3_X1 _34757_ (.A1(_10851_),
    .A2(_10856_),
    .A3(_10876_),
    .ZN(_10892_));
 XNOR2_X1 _34758_ (.A(_10805_),
    .B(_10892_),
    .ZN(_10893_));
 NOR3_X1 _34759_ (.A1(_10883_),
    .A2(_10859_),
    .A3(_10893_),
    .ZN(_10894_));
 NOR2_X1 _34760_ (.A1(_10740_),
    .A2(_10885_),
    .ZN(_10895_));
 AOI21_X1 _34761_ (.A(_10894_),
    .B1(_10895_),
    .B2(_10889_),
    .ZN(_10896_));
 AOI21_X2 _34762_ (.A(_10891_),
    .B1(_10896_),
    .B2(_10869_),
    .ZN(_00011_));
 NOR2_X2 _34763_ (.A1(\g_reduce0[0].adder.b[6] ),
    .A2(_10862_),
    .ZN(_10897_));
 AOI21_X2 _34764_ (.A(net344),
    .B1(_10863_),
    .B2(\g_reduce0[0].adder.a[6] ),
    .ZN(_10898_));
 NAND2_X1 _34765_ (.A1(_10809_),
    .A2(_10807_),
    .ZN(_10899_));
 NOR2_X1 _34766_ (.A1(_10805_),
    .A2(_10857_),
    .ZN(_10900_));
 XNOR2_X2 _34767_ (.A(_10899_),
    .B(_10900_),
    .ZN(_10901_));
 OAI211_X2 _34768_ (.A(_10740_),
    .B(_10901_),
    .C1(_10877_),
    .C2(_10888_),
    .ZN(_10902_));
 OAI21_X1 _34769_ (.A(_10883_),
    .B1(_10859_),
    .B2(_10893_),
    .ZN(_10903_));
 NAND3_X2 _34770_ (.A1(_10231_),
    .A2(_10902_),
    .A3(_10903_),
    .ZN(_10904_));
 AOI21_X4 _34771_ (.A(_10897_),
    .B1(_10898_),
    .B2(_10904_),
    .ZN(_00012_));
 AOI22_X4 _34772_ (.A1(\g_reduce0[0].adder.b[7] ),
    .A2(net344),
    .B1(_10698_),
    .B2(\g_reduce0[0].adder.a[7] ),
    .ZN(_10905_));
 AND3_X1 _34773_ (.A1(_10851_),
    .A2(_10856_),
    .A3(_10876_),
    .ZN(_10906_));
 NAND2_X1 _34774_ (.A1(_10810_),
    .A2(_10906_),
    .ZN(_10907_));
 XOR2_X2 _34775_ (.A(_10835_),
    .B(_10907_),
    .Z(_10908_));
 MUX2_X1 _34776_ (.A(_10908_),
    .B(_10901_),
    .S(_10860_),
    .Z(_10909_));
 OAI21_X2 _34777_ (.A(_10905_),
    .B1(_10909_),
    .B2(_10701_),
    .ZN(_00013_));
 AOI22_X4 _34778_ (.A1(\g_reduce0[0].adder.b[8] ),
    .A2(net344),
    .B1(_10698_),
    .B2(\g_reduce0[0].adder.a[8] ),
    .ZN(_10910_));
 NOR3_X1 _34779_ (.A1(_10836_),
    .A2(_10797_),
    .A3(_10857_),
    .ZN(_10911_));
 NOR2_X1 _34780_ (.A1(_10740_),
    .A2(_10780_),
    .ZN(_10912_));
 OAI21_X1 _34781_ (.A(_10911_),
    .B1(_10912_),
    .B2(_10908_),
    .ZN(_10913_));
 AOI21_X1 _34782_ (.A(_10701_),
    .B1(_10908_),
    .B2(_10883_),
    .ZN(_10914_));
 NAND2_X1 _34783_ (.A1(_10913_),
    .A2(_10914_),
    .ZN(_10915_));
 OR3_X2 _34784_ (.A1(_10786_),
    .A2(_10790_),
    .A3(_10796_),
    .ZN(_10916_));
 NOR2_X1 _34785_ (.A1(_10916_),
    .A2(_10858_),
    .ZN(_10917_));
 AOI21_X1 _34786_ (.A(_10917_),
    .B1(_10911_),
    .B2(_10780_),
    .ZN(_10918_));
 NOR2_X1 _34787_ (.A1(_10883_),
    .A2(_10918_),
    .ZN(_10919_));
 OAI21_X2 _34788_ (.A(_10910_),
    .B1(_10915_),
    .B2(_10919_),
    .ZN(_00014_));
 OAI22_X2 _34789_ (.A1(\g_reduce0[0].adder.b[9] ),
    .A2(_10862_),
    .B1(_10864_),
    .B2(\g_reduce0[0].adder.a[9] ),
    .ZN(_10920_));
 NOR3_X1 _34790_ (.A1(_10883_),
    .A2(_10780_),
    .A3(_10916_),
    .ZN(_10921_));
 NOR3_X1 _34791_ (.A1(_10740_),
    .A2(_10797_),
    .A3(_10858_),
    .ZN(_10922_));
 NAND2_X1 _34792_ (.A1(_10857_),
    .A2(_10892_),
    .ZN(_10923_));
 NOR2_X1 _34793_ (.A1(_10883_),
    .A2(_10836_),
    .ZN(_10924_));
 NAND2_X1 _34794_ (.A1(_10916_),
    .A2(_10892_),
    .ZN(_10925_));
 AOI221_X1 _34795_ (.A(_10780_),
    .B1(_10923_),
    .B2(_10924_),
    .C1(_10925_),
    .C2(_10883_),
    .ZN(_10926_));
 NOR3_X1 _34796_ (.A1(_10740_),
    .A2(_10916_),
    .A3(_10857_),
    .ZN(_10927_));
 AND3_X1 _34797_ (.A1(_10780_),
    .A2(_10916_),
    .A3(_10906_),
    .ZN(_10928_));
 AOI21_X1 _34798_ (.A(_10927_),
    .B1(_10928_),
    .B2(_10740_),
    .ZN(_10929_));
 OAI21_X1 _34799_ (.A(_10869_),
    .B1(_10929_),
    .B2(_10836_),
    .ZN(_10930_));
 NOR4_X1 _34800_ (.A1(_10921_),
    .A2(_10922_),
    .A3(_10926_),
    .A4(_10930_),
    .ZN(_10931_));
 NOR2_X1 _34801_ (.A1(_10920_),
    .A2(_10931_),
    .ZN(_00015_));
 INV_X1 _34802_ (.A(_20478_),
    .ZN(_20484_));
 MUX2_X1 _34803_ (.A(\g_reduce0[0].adder.a[10] ),
    .B(_20483_),
    .S(_10231_),
    .Z(_10932_));
 MUX2_X2 _34804_ (.A(\g_reduce0[0].adder.b[10] ),
    .B(_10932_),
    .S(_10862_),
    .Z(_00001_));
 MUX2_X1 _34805_ (.A(\g_reduce0[0].adder.a[11] ),
    .B(_20491_),
    .S(_10231_),
    .Z(_10933_));
 MUX2_X2 _34806_ (.A(\g_reduce0[0].adder.b[11] ),
    .B(_10933_),
    .S(_10862_),
    .Z(_00002_));
 MUX2_X2 _34807_ (.A(_20356_),
    .B(_00458_),
    .S(_10273_),
    .Z(_10934_));
 NAND2_X1 _34808_ (.A1(_10639_),
    .A2(_20485_),
    .ZN(_10935_));
 XOR2_X1 _34809_ (.A(_10934_),
    .B(_10935_),
    .Z(_10936_));
 XNOR2_X1 _34810_ (.A(_14503_),
    .B(_20495_),
    .ZN(_10937_));
 MUX2_X1 _34811_ (.A(_10936_),
    .B(_10937_),
    .S(_10795_),
    .Z(_10938_));
 XOR2_X1 _34812_ (.A(_20490_),
    .B(_10938_),
    .Z(_10939_));
 MUX2_X1 _34813_ (.A(_10224_),
    .B(_10939_),
    .S(_10231_),
    .Z(_10940_));
 MUX2_X2 _34814_ (.A(\g_reduce0[0].adder.b[12] ),
    .B(_10940_),
    .S(_10862_),
    .Z(_00003_));
 MUX2_X1 _34815_ (.A(_20353_),
    .B(_00461_),
    .S(_10273_),
    .Z(_10941_));
 NOR4_X1 _34816_ (.A1(_10675_),
    .A2(_20478_),
    .A3(_14500_),
    .A4(_10934_),
    .ZN(_10942_));
 XNOR2_X1 _34817_ (.A(_10941_),
    .B(_10942_),
    .ZN(_10943_));
 INV_X1 _34818_ (.A(_20494_),
    .ZN(_10944_));
 INV_X1 _34819_ (.A(_14502_),
    .ZN(_10945_));
 AOI21_X1 _34820_ (.A(_20487_),
    .B1(_20488_),
    .B2(_10945_),
    .ZN(_10946_));
 INV_X1 _34821_ (.A(_20495_),
    .ZN(_10947_));
 OAI21_X1 _34822_ (.A(_10944_),
    .B1(_10946_),
    .B2(_10947_),
    .ZN(_10948_));
 XOR2_X1 _34823_ (.A(_20499_),
    .B(_10948_),
    .Z(_10949_));
 MUX2_X1 _34824_ (.A(_10943_),
    .B(_10949_),
    .S(_10795_),
    .Z(_10950_));
 NOR2_X1 _34825_ (.A1(_10675_),
    .A2(_20486_),
    .ZN(_10951_));
 AOI21_X1 _34826_ (.A(_10951_),
    .B1(_14500_),
    .B2(_10675_),
    .ZN(_10952_));
 NOR2_X1 _34827_ (.A1(_10795_),
    .A2(_10952_),
    .ZN(_10953_));
 AOI21_X2 _34828_ (.A(_10953_),
    .B1(_10795_),
    .B2(_14504_),
    .ZN(_20489_));
 NAND3_X1 _34829_ (.A1(_20482_),
    .A2(_10938_),
    .A3(_20489_),
    .ZN(_10954_));
 XNOR2_X1 _34830_ (.A(_10950_),
    .B(_10954_),
    .ZN(_10955_));
 MUX2_X1 _34831_ (.A(\g_reduce0[0].adder.a[13] ),
    .B(_10955_),
    .S(_10231_),
    .Z(_10956_));
 MUX2_X2 _34832_ (.A(\g_reduce0[0].adder.b[13] ),
    .B(_10956_),
    .S(_10862_),
    .Z(_00004_));
 NOR2_X1 _34833_ (.A1(_10228_),
    .A2(_10362_),
    .ZN(_10957_));
 NOR4_X1 _34834_ (.A1(_10795_),
    .A2(_10934_),
    .A3(_10935_),
    .A4(_10941_),
    .ZN(_10958_));
 OAI21_X1 _34835_ (.A(_10944_),
    .B1(_10947_),
    .B2(_14503_),
    .ZN(_10959_));
 AOI21_X1 _34836_ (.A(_20498_),
    .B1(_10959_),
    .B2(_20499_),
    .ZN(_10960_));
 AOI21_X1 _34837_ (.A(_10958_),
    .B1(_10960_),
    .B2(_10795_),
    .ZN(_10961_));
 NAND3_X1 _34838_ (.A1(_20490_),
    .A2(_10938_),
    .A3(_10950_),
    .ZN(_10962_));
 XNOR2_X1 _34839_ (.A(_10961_),
    .B(_10962_),
    .ZN(_10963_));
 MUX2_X1 _34840_ (.A(_10957_),
    .B(_10362_),
    .S(_10963_),
    .Z(_10964_));
 OAI21_X1 _34841_ (.A(_10225_),
    .B1(_10863_),
    .B2(_10964_),
    .ZN(_10965_));
 AND2_X1 _34842_ (.A1(_10228_),
    .A2(_10292_),
    .ZN(_10966_));
 NOR2_X1 _34843_ (.A1(_10228_),
    .A2(_10700_),
    .ZN(_10967_));
 NOR3_X1 _34844_ (.A1(_10225_),
    .A2(_10966_),
    .A3(_10967_),
    .ZN(_10968_));
 MUX2_X1 _34845_ (.A(_10968_),
    .B(_10966_),
    .S(_10963_),
    .Z(_10969_));
 AOI22_X2 _34846_ (.A1(_10228_),
    .A2(_10227_),
    .B1(_10231_),
    .B2(_10969_),
    .ZN(_10970_));
 NAND2_X2 _34847_ (.A1(_10965_),
    .A2(_10970_),
    .ZN(_00005_));
 OR2_X1 _34848_ (.A1(\g_reduce0[10].adder.a[10] ),
    .A2(\g_reduce0[10].adder.a[13] ),
    .ZN(_10971_));
 OR4_X1 _34849_ (.A1(\g_reduce0[10].adder.a[11] ),
    .A2(\g_reduce0[10].adder.a[12] ),
    .A3(\g_reduce0[10].adder.a[14] ),
    .A4(_10971_),
    .ZN(_10972_));
 CLKBUF_X3 _34850_ (.A(_10972_),
    .Z(_10973_));
 CLKBUF_X2 _34851_ (.A(\g_reduce0[10].adder.b[14] ),
    .Z(_10974_));
 OR2_X1 _34852_ (.A1(\g_reduce0[10].adder.b[10] ),
    .A2(\g_reduce0[10].adder.b[13] ),
    .ZN(_10975_));
 NOR4_X4 _34853_ (.A1(\g_reduce0[10].adder.b[11] ),
    .A2(\g_reduce0[10].adder.b[12] ),
    .A3(_10974_),
    .A4(_10975_),
    .ZN(_10976_));
 INV_X1 _34854_ (.A(_20517_),
    .ZN(_10977_));
 AOI21_X1 _34855_ (.A(_20519_),
    .B1(_20520_),
    .B2(_20522_),
    .ZN(_10978_));
 NOR2_X1 _34856_ (.A1(_10977_),
    .A2(_10978_),
    .ZN(_10979_));
 OAI21_X2 _34857_ (.A(_20514_),
    .B1(_20516_),
    .B2(_10979_),
    .ZN(_10980_));
 INV_X4 _34858_ (.A(_20511_),
    .ZN(_10981_));
 NAND4_X1 _34859_ (.A1(_20514_),
    .A2(_20517_),
    .A3(_20520_),
    .A4(_20523_),
    .ZN(_10982_));
 AOI21_X1 _34860_ (.A(_20525_),
    .B1(_20528_),
    .B2(_20526_),
    .ZN(_10983_));
 NOR2_X1 _34861_ (.A1(_10982_),
    .A2(_10983_),
    .ZN(_10984_));
 CLKBUF_X3 _34862_ (.A(_20544_),
    .Z(_10985_));
 BUF_X4 _34863_ (.A(_20502_),
    .Z(_10986_));
 BUF_X2 _34864_ (.A(_20505_),
    .Z(_10987_));
 INV_X1 _34865_ (.A(_10987_),
    .ZN(_10988_));
 INV_X1 _34866_ (.A(_20508_),
    .ZN(_10989_));
 NOR2_X2 _34867_ (.A1(_10988_),
    .A2(_10989_),
    .ZN(_10990_));
 NAND3_X2 _34868_ (.A1(_10985_),
    .A2(_10986_),
    .A3(_10990_),
    .ZN(_10991_));
 NOR4_X4 _34869_ (.A1(_20513_),
    .A2(_10981_),
    .A3(_10984_),
    .A4(_10991_),
    .ZN(_10992_));
 NAND2_X1 _34870_ (.A1(_20526_),
    .A2(_20529_),
    .ZN(_10993_));
 NOR2_X1 _34871_ (.A1(_10982_),
    .A2(_10993_),
    .ZN(_10994_));
 AND2_X1 _34872_ (.A1(_20532_),
    .A2(_10994_),
    .ZN(_10995_));
 INV_X1 _34873_ (.A(_20535_),
    .ZN(_10996_));
 INV_X1 _34874_ (.A(_20537_),
    .ZN(_10997_));
 INV_X1 _34875_ (.A(\g_reduce0[10].adder.a[0] ),
    .ZN(_10998_));
 OAI21_X1 _34876_ (.A(_20538_),
    .B1(\g_reduce0[10].adder.b[0] ),
    .B2(_10998_),
    .ZN(_10999_));
 AOI21_X1 _34877_ (.A(_10996_),
    .B1(_10997_),
    .B2(_10999_),
    .ZN(_11000_));
 OAI21_X2 _34878_ (.A(_10995_),
    .B1(_11000_),
    .B2(_20534_),
    .ZN(_11001_));
 NAND2_X1 _34879_ (.A1(_20531_),
    .A2(_10994_),
    .ZN(_11002_));
 NAND4_X4 _34880_ (.A1(_10980_),
    .A2(_10992_),
    .A3(_11001_),
    .A4(_11002_),
    .ZN(_11003_));
 INV_X1 _34881_ (.A(_20543_),
    .ZN(_11004_));
 INV_X1 _34882_ (.A(_20504_),
    .ZN(_11005_));
 INV_X1 _34883_ (.A(_20510_),
    .ZN(_11006_));
 AOI21_X1 _34884_ (.A(_20507_),
    .B1(_11006_),
    .B2(_20508_),
    .ZN(_11007_));
 OAI21_X1 _34885_ (.A(_11005_),
    .B1(_11007_),
    .B2(_10988_),
    .ZN(_11008_));
 AOI21_X2 _34886_ (.A(_20501_),
    .B1(_11008_),
    .B2(_10986_),
    .ZN(_11009_));
 INV_X2 _34887_ (.A(_10985_),
    .ZN(_11010_));
 OAI21_X4 _34888_ (.A(_11004_),
    .B1(_11009_),
    .B2(_11010_),
    .ZN(_11011_));
 NAND2_X1 _34889_ (.A1(_11003_),
    .A2(_11011_),
    .ZN(_11012_));
 OAI21_X1 _34890_ (.A(_10973_),
    .B1(_10976_),
    .B2(_11012_),
    .ZN(_11013_));
 MUX2_X1 _34891_ (.A(\g_reduce0[10].adder.a[15] ),
    .B(\g_reduce0[10].adder.b[15] ),
    .S(_11013_),
    .Z(_00022_));
 AND4_X1 _34892_ (.A1(_10980_),
    .A2(_10992_),
    .A3(_11001_),
    .A4(_11002_),
    .ZN(_11014_));
 BUF_X4 _34893_ (.A(_11014_),
    .Z(_11015_));
 INV_X1 _34894_ (.A(_20501_),
    .ZN(_11016_));
 INV_X1 _34895_ (.A(_20507_),
    .ZN(_11017_));
 OAI21_X1 _34896_ (.A(_11017_),
    .B1(_20510_),
    .B2(_10989_),
    .ZN(_11018_));
 AOI21_X1 _34897_ (.A(_20504_),
    .B1(_11018_),
    .B2(_10987_),
    .ZN(_11019_));
 INV_X2 _34898_ (.A(_10986_),
    .ZN(_11020_));
 OAI21_X2 _34899_ (.A(_11016_),
    .B1(_11019_),
    .B2(_11020_),
    .ZN(_11021_));
 AOI21_X4 _34900_ (.A(_20543_),
    .B1(_11021_),
    .B2(_10985_),
    .ZN(_11022_));
 NOR2_X4 _34901_ (.A1(_11015_),
    .A2(_11022_),
    .ZN(_11023_));
 MUX2_X2 _34902_ (.A(\g_reduce0[10].adder.a[10] ),
    .B(\g_reduce0[10].adder.b[10] ),
    .S(_11023_),
    .Z(_20628_));
 NOR2_X1 _34903_ (.A1(\g_reduce0[10].adder.a[12] ),
    .A2(_00472_),
    .ZN(_11024_));
 NOR2_X1 _34904_ (.A1(\g_reduce0[10].adder.a[11] ),
    .A2(_00467_),
    .ZN(_11025_));
 AOI21_X1 _34905_ (.A(_11024_),
    .B1(_11025_),
    .B2(_10987_),
    .ZN(_11026_));
 NAND3_X2 _34906_ (.A1(_11003_),
    .A2(_11011_),
    .A3(_11026_),
    .ZN(_11027_));
 NOR2_X1 _34907_ (.A1(\g_reduce0[10].adder.b[11] ),
    .A2(_20506_),
    .ZN(_11028_));
 NAND2_X1 _34908_ (.A1(_10987_),
    .A2(_11028_),
    .ZN(_11029_));
 OAI221_X2 _34909_ (.A(_11029_),
    .B1(_11022_),
    .B2(_11015_),
    .C1(\g_reduce0[10].adder.b[12] ),
    .C2(_20503_),
    .ZN(_11030_));
 AND3_X1 _34910_ (.A1(_10986_),
    .A2(_11027_),
    .A3(_11030_),
    .ZN(_11031_));
 OR4_X1 _34911_ (.A1(\g_reduce0[10].adder.a[13] ),
    .A2(_00475_),
    .A3(_11015_),
    .A4(_11022_),
    .ZN(_11032_));
 NOR2_X1 _34912_ (.A1(\g_reduce0[10].adder.b[13] ),
    .A2(_20500_),
    .ZN(_11033_));
 OAI21_X1 _34913_ (.A(_11033_),
    .B1(_11022_),
    .B2(_11015_),
    .ZN(_11034_));
 NAND3_X1 _34914_ (.A1(_20540_),
    .A2(_10986_),
    .A3(_10987_),
    .ZN(_11035_));
 NAND3_X2 _34915_ (.A1(_11032_),
    .A2(_11034_),
    .A3(_11035_),
    .ZN(_11036_));
 OAI21_X4 _34916_ (.A(_10985_),
    .B1(_11031_),
    .B2(_11036_),
    .ZN(_11037_));
 NAND3_X2 _34917_ (.A1(_10986_),
    .A2(_11027_),
    .A3(_11030_),
    .ZN(_11038_));
 AND3_X2 _34918_ (.A1(_11032_),
    .A2(_11034_),
    .A3(_11035_),
    .ZN(_11039_));
 NAND3_X4 _34919_ (.A1(_11010_),
    .A2(_11038_),
    .A3(_11039_),
    .ZN(_11040_));
 AND2_X1 _34920_ (.A1(_11027_),
    .A2(_11030_),
    .ZN(_11041_));
 INV_X1 _34921_ (.A(\g_reduce0[10].adder.b[10] ),
    .ZN(_11042_));
 NAND4_X2 _34922_ (.A1(\g_reduce0[10].adder.a[10] ),
    .A2(_11042_),
    .A3(_11003_),
    .A4(_11011_),
    .ZN(_11043_));
 NOR2_X1 _34923_ (.A1(\g_reduce0[10].adder.a[10] ),
    .A2(_11042_),
    .ZN(_11044_));
 OAI21_X1 _34924_ (.A(_11044_),
    .B1(_11022_),
    .B2(_11015_),
    .ZN(_11045_));
 AND3_X1 _34925_ (.A1(_10990_),
    .A2(_11043_),
    .A3(_11045_),
    .ZN(_11046_));
 OAI21_X4 _34926_ (.A(_10986_),
    .B1(_11041_),
    .B2(_11046_),
    .ZN(_11047_));
 NAND2_X2 _34927_ (.A1(_11027_),
    .A2(_11030_),
    .ZN(_11048_));
 NAND3_X2 _34928_ (.A1(_10990_),
    .A2(_11043_),
    .A3(_11045_),
    .ZN(_11049_));
 NAND3_X4 _34929_ (.A1(_11020_),
    .A2(_11048_),
    .A3(_11049_),
    .ZN(_11050_));
 AOI22_X4 _34930_ (.A1(_11037_),
    .A2(_11040_),
    .B1(_11047_),
    .B2(_11050_),
    .ZN(_11051_));
 INV_X1 _34931_ (.A(_20540_),
    .ZN(_11052_));
 OAI21_X1 _34932_ (.A(_11028_),
    .B1(_11022_),
    .B2(_11015_),
    .ZN(_11053_));
 NAND3_X1 _34933_ (.A1(_11003_),
    .A2(_11011_),
    .A3(_11025_),
    .ZN(_11054_));
 AND3_X1 _34934_ (.A1(_11052_),
    .A2(_11053_),
    .A3(_11054_),
    .ZN(_11055_));
 XNOR2_X2 _34935_ (.A(_10987_),
    .B(_11055_),
    .ZN(_11056_));
 CLKBUF_X3 _34936_ (.A(_20541_),
    .Z(_11057_));
 BUF_X4 _34937_ (.A(_11057_),
    .Z(_11058_));
 MUX2_X1 _34938_ (.A(_00470_),
    .B(_20518_),
    .S(_11023_),
    .Z(_11059_));
 CLKBUF_X3 _34939_ (.A(_11023_),
    .Z(_11060_));
 MUX2_X1 _34940_ (.A(_00471_),
    .B(_20521_),
    .S(_11060_),
    .Z(_11061_));
 CLKBUF_X3 _34941_ (.A(_20511_),
    .Z(_11062_));
 BUF_X4 _34942_ (.A(_11062_),
    .Z(_11063_));
 MUX2_X1 _34943_ (.A(_11059_),
    .B(_11061_),
    .S(_11063_),
    .Z(_11064_));
 AND2_X1 _34944_ (.A1(_11058_),
    .A2(_11064_),
    .ZN(_11065_));
 MUX2_X1 _34945_ (.A(_00468_),
    .B(_20524_),
    .S(_11060_),
    .Z(_11066_));
 MUX2_X1 _34946_ (.A(_00469_),
    .B(_20527_),
    .S(_11060_),
    .Z(_11067_));
 MUX2_X1 _34947_ (.A(_11066_),
    .B(_11067_),
    .S(_11063_),
    .Z(_11068_));
 INV_X2 _34948_ (.A(_11057_),
    .ZN(_11069_));
 AOI21_X1 _34949_ (.A(_11065_),
    .B1(_11068_),
    .B2(_11069_),
    .ZN(_11070_));
 NAND2_X1 _34950_ (.A1(_11056_),
    .A2(_11070_),
    .ZN(_11071_));
 MUX2_X1 _34951_ (.A(_00462_),
    .B(_20536_),
    .S(_11060_),
    .Z(_11072_));
 MUX2_X1 _34952_ (.A(_00463_),
    .B(_00464_),
    .S(_11060_),
    .Z(_11073_));
 MUX2_X1 _34953_ (.A(_11072_),
    .B(_11073_),
    .S(_11063_),
    .Z(_11074_));
 NOR2_X1 _34954_ (.A1(_11058_),
    .A2(_11074_),
    .ZN(_11075_));
 AND2_X1 _34955_ (.A1(_20533_),
    .A2(_11060_),
    .ZN(_11076_));
 AOI21_X1 _34956_ (.A(_11076_),
    .B1(_11012_),
    .B2(_00466_),
    .ZN(_11077_));
 NOR2_X1 _34957_ (.A1(_10981_),
    .A2(_11077_),
    .ZN(_11078_));
 MUX2_X1 _34958_ (.A(_00465_),
    .B(_20530_),
    .S(_11060_),
    .Z(_11079_));
 AOI21_X1 _34959_ (.A(_11078_),
    .B1(_11079_),
    .B2(_10981_),
    .ZN(_11080_));
 AOI21_X1 _34960_ (.A(_11075_),
    .B1(_11080_),
    .B2(_11058_),
    .ZN(_11081_));
 OAI21_X1 _34961_ (.A(_11071_),
    .B1(_11081_),
    .B2(_11056_),
    .ZN(_11082_));
 MUX2_X1 _34962_ (.A(_00474_),
    .B(_20515_),
    .S(_11060_),
    .Z(_11083_));
 MUX2_X1 _34963_ (.A(_00473_),
    .B(_20512_),
    .S(_11023_),
    .Z(_11084_));
 MUX2_X1 _34964_ (.A(_11083_),
    .B(_11084_),
    .S(_10981_),
    .Z(_11085_));
 MUX2_X1 _34965_ (.A(_10981_),
    .B(_11085_),
    .S(_11069_),
    .Z(_11086_));
 INV_X1 _34966_ (.A(_11086_),
    .ZN(_11087_));
 NAND2_X1 _34967_ (.A1(_11037_),
    .A2(_11040_),
    .ZN(_11088_));
 NOR3_X2 _34968_ (.A1(_10986_),
    .A2(_11041_),
    .A3(_11046_),
    .ZN(_11089_));
 AOI21_X2 _34969_ (.A(_11020_),
    .B1(_11048_),
    .B2(_11049_),
    .ZN(_11090_));
 NOR2_X2 _34970_ (.A1(_11089_),
    .A2(_11090_),
    .ZN(_11091_));
 XNOR2_X1 _34971_ (.A(_10988_),
    .B(_11055_),
    .ZN(_11092_));
 BUF_X1 _34972_ (.A(_11092_),
    .Z(_11093_));
 AND3_X1 _34973_ (.A1(_11088_),
    .A2(_11091_),
    .A3(_11093_),
    .ZN(_11094_));
 AOI22_X2 _34974_ (.A1(_11051_),
    .A2(_11082_),
    .B1(_11087_),
    .B2(_11094_),
    .ZN(_20608_));
 INV_X1 _34975_ (.A(_20608_),
    .ZN(_20605_));
 AOI21_X4 _34976_ (.A(_11058_),
    .B1(_11084_),
    .B2(_11063_),
    .ZN(_11095_));
 NAND2_X1 _34977_ (.A1(_11062_),
    .A2(_00468_),
    .ZN(_11096_));
 INV_X1 _34978_ (.A(_00471_),
    .ZN(_11097_));
 OAI221_X1 _34979_ (.A(_11096_),
    .B1(_11022_),
    .B2(_11015_),
    .C1(_11063_),
    .C2(_11097_),
    .ZN(_11098_));
 INV_X1 _34980_ (.A(_20524_),
    .ZN(_11099_));
 NAND2_X1 _34981_ (.A1(_11062_),
    .A2(_11099_),
    .ZN(_11100_));
 OAI21_X1 _34982_ (.A(_11100_),
    .B1(_20521_),
    .B2(_11062_),
    .ZN(_11101_));
 NAND3_X1 _34983_ (.A1(_11003_),
    .A2(_11011_),
    .A3(_11101_),
    .ZN(_11102_));
 NAND2_X1 _34984_ (.A1(_11098_),
    .A2(_11102_),
    .ZN(_11103_));
 NOR2_X1 _34985_ (.A1(_11058_),
    .A2(_11103_),
    .ZN(_11104_));
 MUX2_X1 _34986_ (.A(_11059_),
    .B(_11083_),
    .S(_10981_),
    .Z(_11105_));
 AOI21_X1 _34987_ (.A(_11104_),
    .B1(_11105_),
    .B2(_11058_),
    .ZN(_11106_));
 NAND2_X1 _34988_ (.A1(_11062_),
    .A2(_00465_),
    .ZN(_11107_));
 INV_X1 _34989_ (.A(_00469_),
    .ZN(_11108_));
 OAI221_X2 _34990_ (.A(_11107_),
    .B1(_11022_),
    .B2(_11015_),
    .C1(_11063_),
    .C2(_11108_),
    .ZN(_11109_));
 INV_X1 _34991_ (.A(_20530_),
    .ZN(_11110_));
 NAND2_X1 _34992_ (.A1(_11062_),
    .A2(_11110_),
    .ZN(_11111_));
 OAI21_X1 _34993_ (.A(_11111_),
    .B1(_20527_),
    .B2(_11062_),
    .ZN(_11112_));
 NAND3_X1 _34994_ (.A1(_11003_),
    .A2(_11011_),
    .A3(_11112_),
    .ZN(_11113_));
 NAND2_X1 _34995_ (.A1(_11109_),
    .A2(_11113_),
    .ZN(_11114_));
 NAND2_X1 _34996_ (.A1(_11058_),
    .A2(_11114_),
    .ZN(_11115_));
 NOR2_X1 _34997_ (.A1(_10981_),
    .A2(_11072_),
    .ZN(_11116_));
 AOI21_X1 _34998_ (.A(_11116_),
    .B1(_11077_),
    .B2(_10981_),
    .ZN(_11117_));
 OAI21_X1 _34999_ (.A(_11115_),
    .B1(_11117_),
    .B2(_11058_),
    .ZN(_11118_));
 MUX2_X1 _35000_ (.A(_11106_),
    .B(_11118_),
    .S(_11093_),
    .Z(_11119_));
 AOI22_X4 _35001_ (.A1(_11094_),
    .A2(_11095_),
    .B1(_11119_),
    .B2(_11051_),
    .ZN(_14512_));
 INV_X1 _35002_ (.A(_14512_),
    .ZN(_14508_));
 AOI221_X2 _35003_ (.A(_11056_),
    .B1(_11040_),
    .B2(_11037_),
    .C1(_11050_),
    .C2(_11047_),
    .ZN(_11120_));
 BUF_X4 _35004_ (.A(_11120_),
    .Z(_11121_));
 NAND2_X1 _35005_ (.A1(_11095_),
    .A2(_11121_),
    .ZN(_20560_));
 INV_X1 _35006_ (.A(_20560_),
    .ZN(_20564_));
 NAND2_X1 _35007_ (.A1(_11087_),
    .A2(_11121_),
    .ZN(_20553_));
 INV_X1 _35008_ (.A(_20553_),
    .ZN(_20557_));
 NOR2_X1 _35009_ (.A1(_11062_),
    .A2(_11057_),
    .ZN(_11122_));
 MUX2_X1 _35010_ (.A(_00470_),
    .B(_00473_),
    .S(_11057_),
    .Z(_11123_));
 AOI221_X1 _35011_ (.A(_11023_),
    .B1(_11122_),
    .B2(_00474_),
    .C1(_11123_),
    .C2(_11062_),
    .ZN(_11124_));
 MUX2_X1 _35012_ (.A(_20518_),
    .B(_20512_),
    .S(_11057_),
    .Z(_11125_));
 AOI221_X1 _35013_ (.A(_11012_),
    .B1(_11125_),
    .B2(_11062_),
    .C1(_11122_),
    .C2(_20515_),
    .ZN(_11126_));
 OR2_X2 _35014_ (.A1(_11124_),
    .A2(_11126_),
    .ZN(_11127_));
 NAND2_X1 _35015_ (.A1(_11121_),
    .A2(_11127_),
    .ZN(_20589_));
 INV_X1 _35016_ (.A(_20589_),
    .ZN(_20592_));
 NAND2_X2 _35017_ (.A1(_11050_),
    .A2(_11047_),
    .ZN(_11128_));
 NAND2_X1 _35018_ (.A1(_11088_),
    .A2(_11128_),
    .ZN(_11129_));
 NAND2_X4 _35019_ (.A1(_11063_),
    .A2(_11069_),
    .ZN(_11130_));
 MUX2_X1 _35020_ (.A(_11064_),
    .B(_11085_),
    .S(_11058_),
    .Z(_11131_));
 MUX2_X1 _35021_ (.A(_11130_),
    .B(_11131_),
    .S(_11093_),
    .Z(_11132_));
 OR2_X1 _35022_ (.A1(_11129_),
    .A2(_11132_),
    .ZN(_20567_));
 INV_X1 _35023_ (.A(_20567_),
    .ZN(_20571_));
 MUX2_X1 _35024_ (.A(_11095_),
    .B(_11106_),
    .S(_11093_),
    .Z(_11133_));
 AND2_X1 _35025_ (.A1(_11051_),
    .A2(_11133_),
    .ZN(_20575_));
 INV_X1 _35026_ (.A(_20575_),
    .ZN(_20578_));
 NOR2_X1 _35027_ (.A1(_11093_),
    .A2(_11086_),
    .ZN(_11134_));
 AOI21_X1 _35028_ (.A(_11134_),
    .B1(_11070_),
    .B2(_11093_),
    .ZN(_11135_));
 NOR2_X1 _35029_ (.A1(_11129_),
    .A2(_11135_),
    .ZN(_20581_));
 INV_X1 _35030_ (.A(_20581_),
    .ZN(_20585_));
 MUX2_X1 _35031_ (.A(_11103_),
    .B(_11114_),
    .S(_11069_),
    .Z(_11136_));
 MUX2_X1 _35032_ (.A(_11127_),
    .B(_11136_),
    .S(_11093_),
    .Z(_11137_));
 AND2_X1 _35033_ (.A1(_11051_),
    .A2(_11137_),
    .ZN(_20599_));
 INV_X1 _35034_ (.A(_20599_),
    .ZN(_20602_));
 NOR2_X1 _35035_ (.A1(_11069_),
    .A2(_11068_),
    .ZN(_11138_));
 AOI21_X1 _35036_ (.A(_11138_),
    .B1(_11080_),
    .B2(_11069_),
    .ZN(_11139_));
 MUX2_X1 _35037_ (.A(_11131_),
    .B(_11139_),
    .S(_11093_),
    .Z(_11140_));
 NOR2_X1 _35038_ (.A1(_11129_),
    .A2(_11140_),
    .ZN(_11141_));
 NOR2_X4 _35039_ (.A1(_10981_),
    .A2(_11058_),
    .ZN(_11142_));
 AOI21_X2 _35040_ (.A(_11141_),
    .B1(_11142_),
    .B2(_11094_),
    .ZN(_20595_));
 INV_X1 _35041_ (.A(_20595_),
    .ZN(_20550_));
 XOR2_X2 _35042_ (.A(\g_reduce0[10].adder.a[15] ),
    .B(\g_reduce0[10].adder.b[15] ),
    .Z(_11143_));
 BUF_X4 _35043_ (.A(_11143_),
    .Z(_11144_));
 CLKBUF_X2 _35044_ (.A(_20563_),
    .Z(_11145_));
 INV_X2 _35045_ (.A(_11145_),
    .ZN(_11146_));
 INV_X1 _35046_ (.A(_20558_),
    .ZN(_11147_));
 INV_X1 _35047_ (.A(_20591_),
    .ZN(_11148_));
 BUF_X1 _35048_ (.A(_20570_),
    .Z(_11149_));
 INV_X1 _35049_ (.A(_11149_),
    .ZN(_11150_));
 AOI21_X1 _35050_ (.A(_20572_),
    .B1(_20576_),
    .B2(_11150_),
    .ZN(_11151_));
 BUF_X2 _35051_ (.A(_20577_),
    .Z(_11152_));
 BUF_X2 _35052_ (.A(_20584_),
    .Z(_11153_));
 OAI21_X1 _35053_ (.A(_11152_),
    .B1(_11153_),
    .B2(_20583_),
    .ZN(_11154_));
 INV_X1 _35054_ (.A(_11154_),
    .ZN(_11155_));
 NAND2_X1 _35055_ (.A1(_11150_),
    .A2(_11155_),
    .ZN(_11156_));
 OR2_X1 _35056_ (.A1(_20583_),
    .A2(_20600_),
    .ZN(_11157_));
 INV_X1 _35057_ (.A(_20551_),
    .ZN(_11158_));
 INV_X1 _35058_ (.A(_20552_),
    .ZN(_11159_));
 AOI21_X1 _35059_ (.A(_20545_),
    .B1(_14507_),
    .B2(_20546_),
    .ZN(_11160_));
 OAI21_X2 _35060_ (.A(_11158_),
    .B1(_11159_),
    .B2(_11160_),
    .ZN(_11161_));
 BUF_X2 _35061_ (.A(_20601_),
    .Z(_11162_));
 AOI21_X1 _35062_ (.A(_11157_),
    .B1(_11161_),
    .B2(_11162_),
    .ZN(_11163_));
 OAI21_X1 _35063_ (.A(_11151_),
    .B1(_11156_),
    .B2(_11163_),
    .ZN(_11164_));
 AOI21_X1 _35064_ (.A(_20593_),
    .B1(_11148_),
    .B2(_11164_),
    .ZN(_11165_));
 BUF_X2 _35065_ (.A(_20556_),
    .Z(_11166_));
 OAI21_X2 _35066_ (.A(_11147_),
    .B1(_11165_),
    .B2(_11166_),
    .ZN(_11167_));
 AOI21_X4 _35067_ (.A(_20565_),
    .B1(_11146_),
    .B2(_11167_),
    .ZN(_11168_));
 NOR2_X2 _35068_ (.A1(_11144_),
    .A2(_11168_),
    .ZN(_11169_));
 XNOR2_X2 _35069_ (.A(\g_reduce0[10].adder.a[15] ),
    .B(\g_reduce0[10].adder.b[15] ),
    .ZN(_11170_));
 BUF_X4 _35070_ (.A(_11170_),
    .Z(_11171_));
 INV_X1 _35071_ (.A(_20590_),
    .ZN(_11172_));
 OAI21_X1 _35072_ (.A(_20591_),
    .B1(_20569_),
    .B2(_11149_),
    .ZN(_11173_));
 NAND2_X1 _35073_ (.A1(_11172_),
    .A2(_11173_),
    .ZN(_11174_));
 NOR2_X1 _35074_ (.A1(_20590_),
    .A2(_20569_),
    .ZN(_11175_));
 INV_X1 _35075_ (.A(_20579_),
    .ZN(_11176_));
 INV_X1 _35076_ (.A(_20586_),
    .ZN(_11177_));
 INV_X1 _35077_ (.A(_20603_),
    .ZN(_11178_));
 NAND3_X1 _35078_ (.A1(_11176_),
    .A2(_11177_),
    .A3(_11178_),
    .ZN(_11179_));
 INV_X1 _35079_ (.A(_20596_),
    .ZN(_11180_));
 INV_X1 _35080_ (.A(_20597_),
    .ZN(_11181_));
 AOI21_X1 _35081_ (.A(_20547_),
    .B1(_14513_),
    .B2(_20548_),
    .ZN(_11182_));
 OAI21_X1 _35082_ (.A(_11180_),
    .B1(_11181_),
    .B2(_11182_),
    .ZN(_11183_));
 INV_X1 _35083_ (.A(_11162_),
    .ZN(_11184_));
 AOI21_X1 _35084_ (.A(_11179_),
    .B1(_11183_),
    .B2(_11184_),
    .ZN(_11185_));
 AOI21_X1 _35085_ (.A(_11152_),
    .B1(_11153_),
    .B2(_11177_),
    .ZN(_11186_));
 NOR2_X1 _35086_ (.A1(_20579_),
    .A2(_11186_),
    .ZN(_11187_));
 OAI21_X1 _35087_ (.A(_11175_),
    .B1(_11185_),
    .B2(_11187_),
    .ZN(_11188_));
 AND3_X1 _35088_ (.A1(_11166_),
    .A2(_11174_),
    .A3(_11188_),
    .ZN(_11189_));
 OAI21_X1 _35089_ (.A(_11145_),
    .B1(_20555_),
    .B2(_11189_),
    .ZN(_11190_));
 INV_X1 _35090_ (.A(_20562_),
    .ZN(_11191_));
 AOI21_X2 _35091_ (.A(_11171_),
    .B1(_11190_),
    .B2(_11191_),
    .ZN(_11192_));
 NOR2_X1 _35092_ (.A1(_11130_),
    .A2(_11192_),
    .ZN(_11193_));
 AOI21_X4 _35093_ (.A(_11169_),
    .B1(_11193_),
    .B2(_11121_),
    .ZN(_11194_));
 AOI21_X1 _35094_ (.A(_20596_),
    .B1(_14514_),
    .B2(_20597_),
    .ZN(_11195_));
 OAI21_X1 _35095_ (.A(_11178_),
    .B1(_11195_),
    .B2(_11162_),
    .ZN(_11196_));
 INV_X1 _35096_ (.A(_11153_),
    .ZN(_11197_));
 AOI21_X2 _35097_ (.A(_20586_),
    .B1(_11196_),
    .B2(_11197_),
    .ZN(_11198_));
 OAI211_X2 _35098_ (.A(_11176_),
    .B(_11175_),
    .C1(_11198_),
    .C2(_11152_),
    .ZN(_11199_));
 AND3_X1 _35099_ (.A1(_11166_),
    .A2(_11174_),
    .A3(_11199_),
    .ZN(_11200_));
 OR2_X1 _35100_ (.A1(_20555_),
    .A2(_11170_),
    .ZN(_11201_));
 NOR3_X1 _35101_ (.A1(_20562_),
    .A2(_11200_),
    .A3(_11201_),
    .ZN(_11202_));
 MUX2_X1 _35102_ (.A(_20558_),
    .B(_11191_),
    .S(_11144_),
    .Z(_11203_));
 INV_X1 _35103_ (.A(_20572_),
    .ZN(_11204_));
 NOR2_X1 _35104_ (.A1(_20583_),
    .A2(_20600_),
    .ZN(_11205_));
 AOI21_X1 _35105_ (.A(_20551_),
    .B1(_14510_),
    .B2(_20552_),
    .ZN(_11206_));
 OAI21_X1 _35106_ (.A(_11205_),
    .B1(_11206_),
    .B2(_11184_),
    .ZN(_11207_));
 AOI21_X1 _35107_ (.A(_20576_),
    .B1(_11155_),
    .B2(_11207_),
    .ZN(_11208_));
 OAI21_X1 _35108_ (.A(_11204_),
    .B1(_11208_),
    .B2(_11149_),
    .ZN(_11209_));
 AOI21_X1 _35109_ (.A(_20593_),
    .B1(_11148_),
    .B2(_11209_),
    .ZN(_11210_));
 NOR3_X1 _35110_ (.A1(_11166_),
    .A2(_11145_),
    .A3(_11210_),
    .ZN(_11211_));
 OR2_X1 _35111_ (.A1(_20565_),
    .A2(_11211_),
    .ZN(_11212_));
 AOI221_X2 _35112_ (.A(_11202_),
    .B1(_11203_),
    .B2(_11146_),
    .C1(_11212_),
    .C2(_11171_),
    .ZN(_11213_));
 INV_X2 _35113_ (.A(_11213_),
    .ZN(_11214_));
 NAND3_X2 _35114_ (.A1(_11121_),
    .A2(_11142_),
    .A3(_11214_),
    .ZN(_11215_));
 NOR3_X2 _35115_ (.A1(_10985_),
    .A2(_11031_),
    .A3(_11036_),
    .ZN(_11216_));
 AOI21_X2 _35116_ (.A(_11010_),
    .B1(_11038_),
    .B2(_11039_),
    .ZN(_11217_));
 OAI221_X2 _35117_ (.A(_11093_),
    .B1(_11216_),
    .B2(_11217_),
    .C1(_11089_),
    .C2(_11090_),
    .ZN(_11218_));
 OAI21_X2 _35118_ (.A(_11213_),
    .B1(_11130_),
    .B2(_11218_),
    .ZN(_11219_));
 NAND2_X4 _35119_ (.A1(_11215_),
    .A2(_11219_),
    .ZN(_11220_));
 AND2_X1 _35120_ (.A1(_11147_),
    .A2(_11165_),
    .ZN(_11221_));
 INV_X1 _35121_ (.A(_11166_),
    .ZN(_11222_));
 OAI21_X2 _35122_ (.A(_11171_),
    .B1(_20558_),
    .B2(_11222_),
    .ZN(_11223_));
 OAI22_X4 _35123_ (.A1(_11189_),
    .A2(_11201_),
    .B1(_11221_),
    .B2(_11223_),
    .ZN(_11224_));
 XNOR2_X2 _35124_ (.A(_11146_),
    .B(_11224_),
    .ZN(_11225_));
 AND2_X1 _35125_ (.A1(_11174_),
    .A2(_11199_),
    .ZN(_11226_));
 MUX2_X1 _35126_ (.A(_11210_),
    .B(_11226_),
    .S(_11143_),
    .Z(_11227_));
 XNOR2_X2 _35127_ (.A(_11166_),
    .B(_11227_),
    .ZN(_11228_));
 NOR3_X1 _35128_ (.A1(_11150_),
    .A2(_11187_),
    .A3(_11185_),
    .ZN(_11229_));
 NOR2_X1 _35129_ (.A1(_20569_),
    .A2(_11229_),
    .ZN(_11230_));
 MUX2_X1 _35130_ (.A(_11164_),
    .B(_11230_),
    .S(_11144_),
    .Z(_11231_));
 XNOR2_X2 _35131_ (.A(_20591_),
    .B(_11231_),
    .ZN(_11232_));
 OAI21_X1 _35132_ (.A(_11176_),
    .B1(_11152_),
    .B2(_11198_),
    .ZN(_11233_));
 MUX2_X1 _35133_ (.A(_11233_),
    .B(_11208_),
    .S(_11170_),
    .Z(_11234_));
 XNOR2_X2 _35134_ (.A(_11149_),
    .B(_11234_),
    .ZN(_11235_));
 AOI21_X1 _35135_ (.A(_20603_),
    .B1(_11183_),
    .B2(_11184_),
    .ZN(_11236_));
 OAI21_X1 _35136_ (.A(_11177_),
    .B1(_11236_),
    .B2(_11153_),
    .ZN(_11237_));
 AOI21_X1 _35137_ (.A(_20600_),
    .B1(_11161_),
    .B2(_11162_),
    .ZN(_11238_));
 OR2_X1 _35138_ (.A1(_11197_),
    .A2(_11238_),
    .ZN(_11239_));
 NOR2_X1 _35139_ (.A1(_20583_),
    .A2(_11143_),
    .ZN(_11240_));
 AOI22_X2 _35140_ (.A1(_11144_),
    .A2(_11237_),
    .B1(_11239_),
    .B2(_11240_),
    .ZN(_11241_));
 XOR2_X2 _35141_ (.A(_11152_),
    .B(_11241_),
    .Z(_11242_));
 AND2_X1 _35142_ (.A1(_11235_),
    .A2(_11242_),
    .ZN(_11243_));
 OAI21_X1 _35143_ (.A(_11228_),
    .B1(_11232_),
    .B2(_11243_),
    .ZN(_11244_));
 NAND2_X2 _35144_ (.A1(_11225_),
    .A2(_11244_),
    .ZN(_11245_));
 NAND2_X4 _35145_ (.A1(_11228_),
    .A2(_11235_),
    .ZN(_11246_));
 INV_X1 _35146_ (.A(_11206_),
    .ZN(_11247_));
 AOI21_X1 _35147_ (.A(_20600_),
    .B1(_11247_),
    .B2(_11162_),
    .ZN(_11248_));
 MUX2_X2 _35148_ (.A(_11196_),
    .B(_11248_),
    .S(_11170_),
    .Z(_11249_));
 XNOR2_X2 _35149_ (.A(_11153_),
    .B(_11249_),
    .ZN(_11250_));
 NOR2_X1 _35150_ (.A1(_11170_),
    .A2(_11183_),
    .ZN(_11251_));
 AOI21_X2 _35151_ (.A(_11251_),
    .B1(_11161_),
    .B2(_11170_),
    .ZN(_11252_));
 XNOR2_X2 _35152_ (.A(_11162_),
    .B(_11252_),
    .ZN(_11253_));
 XOR2_X1 _35153_ (.A(_14510_),
    .B(_20552_),
    .Z(_11254_));
 NAND2_X1 _35154_ (.A1(_11171_),
    .A2(_11254_),
    .ZN(_11255_));
 XOR2_X1 _35155_ (.A(_14514_),
    .B(_20597_),
    .Z(_11256_));
 NAND2_X1 _35156_ (.A1(_11144_),
    .A2(_11256_),
    .ZN(_11257_));
 AND2_X2 _35157_ (.A1(_11255_),
    .A2(_11257_),
    .ZN(_11258_));
 INV_X1 _35158_ (.A(_14515_),
    .ZN(_11259_));
 INV_X1 _35159_ (.A(_14511_),
    .ZN(_11260_));
 MUX2_X2 _35160_ (.A(_11259_),
    .B(_11260_),
    .S(_11171_),
    .Z(_11261_));
 AOI21_X1 _35161_ (.A(_11253_),
    .B1(_11258_),
    .B2(_11261_),
    .ZN(_11262_));
 NOR3_X2 _35162_ (.A1(_11246_),
    .A2(_11250_),
    .A3(_11262_),
    .ZN(_11263_));
 OR2_X1 _35163_ (.A1(_11245_),
    .A2(_11263_),
    .ZN(_11264_));
 AND4_X2 _35164_ (.A1(_11050_),
    .A2(_11047_),
    .A3(_11092_),
    .A4(_11127_),
    .ZN(_11265_));
 XNOR2_X2 _35165_ (.A(_11197_),
    .B(_11249_),
    .ZN(_11266_));
 NAND2_X2 _35166_ (.A1(_11266_),
    .A2(_11258_),
    .ZN(_11267_));
 OR2_X1 _35167_ (.A1(_20609_),
    .A2(_11171_),
    .ZN(_11268_));
 OR3_X1 _35168_ (.A1(_11246_),
    .A2(_11267_),
    .A3(_11268_),
    .ZN(_11269_));
 NAND2_X1 _35169_ (.A1(_11063_),
    .A2(_11057_),
    .ZN(_11270_));
 MUX2_X1 _35170_ (.A(_00464_),
    .B(_20533_),
    .S(_11057_),
    .Z(_11271_));
 OAI221_X1 _35171_ (.A(_11023_),
    .B1(_11270_),
    .B2(_20536_),
    .C1(_11271_),
    .C2(_11063_),
    .ZN(_11272_));
 MUX2_X1 _35172_ (.A(_00463_),
    .B(_00466_),
    .S(_11057_),
    .Z(_11273_));
 OAI221_X2 _35173_ (.A(_11012_),
    .B1(_11270_),
    .B2(_00462_),
    .C1(_11273_),
    .C2(_11063_),
    .ZN(_11274_));
 AND2_X1 _35174_ (.A1(_11272_),
    .A2(_11274_),
    .ZN(_11275_));
 MUX2_X2 _35175_ (.A(_11136_),
    .B(_11275_),
    .S(_11092_),
    .Z(_11276_));
 AOI211_X2 _35176_ (.A(_11265_),
    .B(_11269_),
    .C1(_11128_),
    .C2(_11276_),
    .ZN(_11277_));
 OR2_X1 _35177_ (.A1(_11246_),
    .A2(_11267_),
    .ZN(_11278_));
 OR3_X1 _35178_ (.A1(_11217_),
    .A2(_11216_),
    .A3(_11268_),
    .ZN(_11279_));
 NOR2_X1 _35179_ (.A1(_20607_),
    .A2(_11144_),
    .ZN(_11280_));
 OAI21_X1 _35180_ (.A(_11280_),
    .B1(_11216_),
    .B2(_11217_),
    .ZN(_11281_));
 AOI21_X2 _35181_ (.A(_11278_),
    .B1(_11279_),
    .B2(_11281_),
    .ZN(_11282_));
 NAND4_X2 _35182_ (.A1(_11050_),
    .A2(_11047_),
    .A3(_11093_),
    .A4(_11127_),
    .ZN(_11283_));
 AND2_X1 _35183_ (.A1(_11098_),
    .A2(_11102_),
    .ZN(_11284_));
 AND2_X1 _35184_ (.A1(_11109_),
    .A2(_11113_),
    .ZN(_11285_));
 MUX2_X1 _35185_ (.A(_11284_),
    .B(_11285_),
    .S(_11069_),
    .Z(_11286_));
 NAND2_X1 _35186_ (.A1(_11272_),
    .A2(_11274_),
    .ZN(_11287_));
 MUX2_X1 _35187_ (.A(_11286_),
    .B(_11287_),
    .S(_11092_),
    .Z(_11288_));
 OAI21_X2 _35188_ (.A(_11283_),
    .B1(_11288_),
    .B2(_11091_),
    .ZN(_11289_));
 AOI211_X2 _35189_ (.A(_11264_),
    .B(_11277_),
    .C1(_11282_),
    .C2(_11289_),
    .ZN(_11290_));
 OAI21_X1 _35190_ (.A(_11194_),
    .B1(_11220_),
    .B2(_11290_),
    .ZN(_20611_));
 INV_X2 _35191_ (.A(_20611_),
    .ZN(_20613_));
 BUF_X2 _35192_ (.A(_20616_),
    .Z(_11291_));
 OR2_X1 _35193_ (.A1(_11130_),
    .A2(_11192_),
    .ZN(_11292_));
 OAI22_X4 _35194_ (.A1(_11218_),
    .A2(_11292_),
    .B1(_11168_),
    .B2(_11144_),
    .ZN(_11293_));
 NOR3_X4 _35195_ (.A1(_11218_),
    .A2(_11130_),
    .A3(_11213_),
    .ZN(_11294_));
 AOI21_X4 _35196_ (.A(_11214_),
    .B1(_11142_),
    .B2(_11121_),
    .ZN(_11295_));
 XNOR2_X2 _35197_ (.A(_11145_),
    .B(_11224_),
    .ZN(_11296_));
 OR3_X4 _35198_ (.A1(_11296_),
    .A2(_11232_),
    .A3(_11246_),
    .ZN(_11297_));
 NOR3_X4 _35199_ (.A1(_11242_),
    .A2(_11253_),
    .A3(_11267_),
    .ZN(_11298_));
 NOR2_X4 _35200_ (.A1(_11297_),
    .A2(_11298_),
    .ZN(_11299_));
 NOR4_X4 _35201_ (.A1(_11293_),
    .A2(_11294_),
    .A3(_11295_),
    .A4(_11299_),
    .ZN(_11300_));
 XNOR2_X2 _35202_ (.A(_11291_),
    .B(_11300_),
    .ZN(_11301_));
 INV_X4 _35203_ (.A(_11301_),
    .ZN(_20636_));
 AND4_X2 _35204_ (.A1(_11121_),
    .A2(_11142_),
    .A3(_11192_),
    .A4(_11213_),
    .ZN(_11302_));
 OR2_X1 _35205_ (.A1(_11169_),
    .A2(_11213_),
    .ZN(_11303_));
 AOI21_X4 _35206_ (.A(_11303_),
    .B1(_11142_),
    .B2(_11121_),
    .ZN(_11304_));
 NOR2_X4 _35207_ (.A1(_11302_),
    .A2(_11304_),
    .ZN(_11305_));
 CLKBUF_X3 _35208_ (.A(_11305_),
    .Z(_11306_));
 CLKBUF_X3 _35209_ (.A(_20612_),
    .Z(_11307_));
 BUF_X2 _35210_ (.A(_11307_),
    .Z(_11308_));
 NAND2_X1 _35211_ (.A1(_11308_),
    .A2(_11261_),
    .ZN(_11309_));
 AND2_X1 _35212_ (.A1(_20607_),
    .A2(_11171_),
    .ZN(_11310_));
 AOI21_X4 _35213_ (.A(_11310_),
    .B1(_11144_),
    .B2(_20609_),
    .ZN(_11311_));
 OAI21_X1 _35214_ (.A(_11309_),
    .B1(_11311_),
    .B2(_11308_),
    .ZN(_11312_));
 NAND2_X1 _35215_ (.A1(_11306_),
    .A2(_11312_),
    .ZN(_11313_));
 NOR2_X4 _35216_ (.A1(_11293_),
    .A2(_11220_),
    .ZN(_11314_));
 NOR3_X2 _35217_ (.A1(_11296_),
    .A2(_11232_),
    .A3(_11246_),
    .ZN(_11315_));
 NOR2_X1 _35218_ (.A1(_11291_),
    .A2(_11315_),
    .ZN(_11316_));
 NAND2_X1 _35219_ (.A1(_11291_),
    .A2(_11299_),
    .ZN(_11317_));
 NAND2_X1 _35220_ (.A1(_11225_),
    .A2(_11228_),
    .ZN(_11318_));
 NAND2_X1 _35221_ (.A1(_11255_),
    .A2(_11257_),
    .ZN(_11319_));
 NOR3_X1 _35222_ (.A1(_11260_),
    .A2(_20607_),
    .A3(_11144_),
    .ZN(_11320_));
 NOR3_X1 _35223_ (.A1(_11259_),
    .A2(_20609_),
    .A3(_11171_),
    .ZN(_11321_));
 NOR4_X1 _35224_ (.A1(_11253_),
    .A2(_11319_),
    .A3(_11320_),
    .A4(_11321_),
    .ZN(_11322_));
 NOR3_X1 _35225_ (.A1(_11242_),
    .A2(_11250_),
    .A3(_11322_),
    .ZN(_11323_));
 NOR2_X1 _35226_ (.A1(_11232_),
    .A2(_11323_),
    .ZN(_11324_));
 AOI21_X4 _35227_ (.A(_11318_),
    .B1(_11324_),
    .B2(_11235_),
    .ZN(_11325_));
 AOI21_X2 _35228_ (.A(_11317_),
    .B1(_11325_),
    .B2(_11290_),
    .ZN(_11326_));
 OAI21_X4 _35229_ (.A(_11314_),
    .B1(_11316_),
    .B2(_11326_),
    .ZN(_11327_));
 BUF_X2 _35230_ (.A(_14517_),
    .Z(_11328_));
 INV_X2 _35231_ (.A(_11328_),
    .ZN(_11329_));
 BUF_X4 _35232_ (.A(_11329_),
    .Z(_11330_));
 CLKBUF_X3 _35233_ (.A(_11290_),
    .Z(_11331_));
 AOI22_X2 _35234_ (.A1(_11051_),
    .A2(_11276_),
    .B1(_11265_),
    .B2(_11088_),
    .ZN(_11332_));
 XNOR2_X2 _35235_ (.A(_11171_),
    .B(_11332_),
    .ZN(_11333_));
 NOR3_X2 _35236_ (.A1(_11330_),
    .A2(_11331_),
    .A3(_11333_),
    .ZN(_11334_));
 NAND2_X1 _35237_ (.A1(_11328_),
    .A2(_11311_),
    .ZN(_11335_));
 AOI21_X1 _35238_ (.A(_11334_),
    .B1(_11335_),
    .B2(_20613_),
    .ZN(_11336_));
 OAI21_X1 _35239_ (.A(_11313_),
    .B1(_11327_),
    .B2(_11336_),
    .ZN(_11337_));
 CLKBUF_X3 _35240_ (.A(_11328_),
    .Z(_11338_));
 OAI21_X2 _35241_ (.A(_11333_),
    .B1(_11290_),
    .B2(_11220_),
    .ZN(_11339_));
 NAND3_X2 _35242_ (.A1(_11338_),
    .A2(_11194_),
    .A3(_11339_),
    .ZN(_11340_));
 MUX2_X1 _35243_ (.A(_11333_),
    .B(_11311_),
    .S(_11307_),
    .Z(_11341_));
 OAI22_X4 _35244_ (.A1(_11327_),
    .A2(_11340_),
    .B1(_11341_),
    .B2(_11314_),
    .ZN(_11342_));
 AND2_X1 _35245_ (.A1(_11337_),
    .A2(_11342_),
    .ZN(_20619_));
 NOR4_X4 _35246_ (.A1(\g_reduce0[10].adder.a[11] ),
    .A2(\g_reduce0[10].adder.a[12] ),
    .A3(\g_reduce0[10].adder.a[14] ),
    .A4(_10971_),
    .ZN(_11343_));
 OR4_X1 _35247_ (.A1(\g_reduce0[10].adder.b[11] ),
    .A2(\g_reduce0[10].adder.b[12] ),
    .A3(_10974_),
    .A4(_10975_),
    .ZN(_11344_));
 BUF_X2 _35248_ (.A(_11344_),
    .Z(_11345_));
 NOR2_X1 _35249_ (.A1(_11343_),
    .A2(_11345_),
    .ZN(_11346_));
 AOI22_X1 _35250_ (.A1(\g_reduce0[10].adder.b[0] ),
    .A2(_11343_),
    .B1(_11346_),
    .B2(\g_reduce0[10].adder.a[0] ),
    .ZN(_11347_));
 INV_X1 _35251_ (.A(_20621_),
    .ZN(_11348_));
 NOR2_X1 _35252_ (.A1(_11327_),
    .A2(_11336_),
    .ZN(_11349_));
 AOI21_X1 _35253_ (.A(_11349_),
    .B1(_11312_),
    .B2(_11306_),
    .ZN(_11350_));
 INV_X1 _35254_ (.A(_11325_),
    .ZN(_11351_));
 NOR2_X1 _35255_ (.A1(_11245_),
    .A2(_11263_),
    .ZN(_11352_));
 NOR3_X1 _35256_ (.A1(_11246_),
    .A2(_11267_),
    .A3(_11268_),
    .ZN(_11353_));
 OAI211_X2 _35257_ (.A(_11283_),
    .B(_11353_),
    .C1(_11091_),
    .C2(_11288_),
    .ZN(_11354_));
 NOR2_X1 _35258_ (.A1(_11246_),
    .A2(_11267_),
    .ZN(_11355_));
 NOR3_X1 _35259_ (.A1(_11217_),
    .A2(_11216_),
    .A3(_11268_),
    .ZN(_11356_));
 OR2_X1 _35260_ (.A1(_20607_),
    .A2(_11144_),
    .ZN(_11357_));
 AOI21_X1 _35261_ (.A(_11357_),
    .B1(_11040_),
    .B2(_11037_),
    .ZN(_11358_));
 OAI21_X2 _35262_ (.A(_11355_),
    .B1(_11356_),
    .B2(_11358_),
    .ZN(_11359_));
 AOI21_X2 _35263_ (.A(_11265_),
    .B1(_11276_),
    .B2(_11128_),
    .ZN(_11360_));
 OAI211_X4 _35264_ (.A(_11352_),
    .B(_11354_),
    .C1(_11359_),
    .C2(_11360_),
    .ZN(_11361_));
 OAI21_X2 _35265_ (.A(_11299_),
    .B1(_11351_),
    .B2(_11361_),
    .ZN(_11362_));
 NOR2_X2 _35266_ (.A1(_11297_),
    .A2(_11305_),
    .ZN(_11363_));
 AOI21_X4 _35267_ (.A(_11293_),
    .B1(_11362_),
    .B2(_11363_),
    .ZN(_20641_));
 AND3_X1 _35268_ (.A1(_20614_),
    .A2(_20636_),
    .A3(_20641_),
    .ZN(_11364_));
 OAI21_X1 _35269_ (.A(_11350_),
    .B1(_11364_),
    .B2(_11306_),
    .ZN(_11365_));
 MUX2_X1 _35270_ (.A(_11350_),
    .B(_11365_),
    .S(_11342_),
    .Z(_11366_));
 CLKBUF_X3 _35271_ (.A(_11308_),
    .Z(_11367_));
 CLKBUF_X3 _35272_ (.A(_11194_),
    .Z(_11368_));
 OR2_X1 _35273_ (.A1(_11367_),
    .A2(_11368_),
    .ZN(_11369_));
 NOR2_X1 _35274_ (.A1(_11294_),
    .A2(_11295_),
    .ZN(_11370_));
 CLKBUF_X3 _35275_ (.A(_11370_),
    .Z(_11371_));
 NAND2_X1 _35276_ (.A1(_11371_),
    .A2(_11228_),
    .ZN(_11372_));
 NAND2_X1 _35277_ (.A1(_11368_),
    .A2(_11372_),
    .ZN(_11373_));
 AOI211_X2 _35278_ (.A(_11263_),
    .B(_11277_),
    .C1(_11282_),
    .C2(_11289_),
    .ZN(_11374_));
 CLKBUF_X3 _35279_ (.A(_11220_),
    .Z(_11375_));
 OAI21_X1 _35280_ (.A(_11225_),
    .B1(_11374_),
    .B2(_11375_),
    .ZN(_11376_));
 NAND2_X1 _35281_ (.A1(_11330_),
    .A2(_11376_),
    .ZN(_11377_));
 MUX2_X1 _35282_ (.A(_11253_),
    .B(_11261_),
    .S(_11329_),
    .Z(_11378_));
 AND2_X1 _35283_ (.A1(_11225_),
    .A2(_11244_),
    .ZN(_11379_));
 NOR2_X1 _35284_ (.A1(_11328_),
    .A2(_11311_),
    .ZN(_11380_));
 AOI21_X1 _35285_ (.A(_11380_),
    .B1(_11319_),
    .B2(_11328_),
    .ZN(_11381_));
 NOR2_X1 _35286_ (.A1(_11379_),
    .A2(_11381_),
    .ZN(_11382_));
 MUX2_X1 _35287_ (.A(_11378_),
    .B(_11382_),
    .S(_11371_),
    .Z(_11383_));
 NOR3_X1 _35288_ (.A1(_11294_),
    .A2(_11295_),
    .A3(_11381_),
    .ZN(_11384_));
 MUX2_X1 _35289_ (.A(_14515_),
    .B(_14511_),
    .S(_11171_),
    .Z(_11385_));
 NAND2_X1 _35290_ (.A1(_11329_),
    .A2(_11385_),
    .ZN(_11386_));
 OAI21_X1 _35291_ (.A(_11386_),
    .B1(_11253_),
    .B2(_11329_),
    .ZN(_11387_));
 NOR2_X1 _35292_ (.A1(_11245_),
    .A2(_11387_),
    .ZN(_11388_));
 MUX2_X1 _35293_ (.A(_11384_),
    .B(_11388_),
    .S(_11374_),
    .Z(_11389_));
 OAI21_X2 _35294_ (.A(_11194_),
    .B1(_11383_),
    .B2(_11389_),
    .ZN(_11390_));
 OAI22_X1 _35295_ (.A1(_11373_),
    .A2(_11377_),
    .B1(_11390_),
    .B2(_20641_),
    .ZN(_11391_));
 NOR2_X4 _35296_ (.A1(_11305_),
    .A2(_11301_),
    .ZN(_11392_));
 NAND2_X1 _35297_ (.A1(_11391_),
    .A2(_11392_),
    .ZN(_11393_));
 NOR3_X1 _35298_ (.A1(_11294_),
    .A2(_11295_),
    .A3(_11250_),
    .ZN(_11394_));
 AOI21_X1 _35299_ (.A(_11293_),
    .B1(_11361_),
    .B2(_11394_),
    .ZN(_11395_));
 NOR2_X1 _35300_ (.A1(_11375_),
    .A2(_11331_),
    .ZN(_11396_));
 OAI21_X2 _35301_ (.A(_11395_),
    .B1(_11396_),
    .B2(_11242_),
    .ZN(_11397_));
 NOR2_X1 _35302_ (.A1(_11296_),
    .A2(_11228_),
    .ZN(_11398_));
 NOR3_X1 _35303_ (.A1(_11294_),
    .A2(_11295_),
    .A3(_11398_),
    .ZN(_11399_));
 XNOR2_X1 _35304_ (.A(_11148_),
    .B(_11231_),
    .ZN(_11400_));
 OAI33_X1 _35305_ (.A1(_11235_),
    .A2(_11379_),
    .A3(_11306_),
    .B1(_11399_),
    .B2(_11293_),
    .B3(_11400_),
    .ZN(_11401_));
 NOR2_X1 _35306_ (.A1(_11330_),
    .A2(_11401_),
    .ZN(_11402_));
 NAND4_X2 _35307_ (.A1(_11368_),
    .A2(_11339_),
    .A3(_11362_),
    .A4(_11363_),
    .ZN(_11403_));
 AOI22_X4 _35308_ (.A1(_11330_),
    .A2(_11397_),
    .B1(_11402_),
    .B2(_11403_),
    .ZN(_11404_));
 NOR2_X1 _35309_ (.A1(_11305_),
    .A2(_20636_),
    .ZN(_11405_));
 NAND2_X1 _35310_ (.A1(_11404_),
    .A2(_11405_),
    .ZN(_11406_));
 AND3_X2 _35311_ (.A1(_11369_),
    .A2(_11393_),
    .A3(_11406_),
    .ZN(_11407_));
 OAI21_X1 _35312_ (.A(_11311_),
    .B1(_11331_),
    .B2(_11220_),
    .ZN(_11408_));
 NAND3_X1 _35313_ (.A1(_11371_),
    .A2(_11361_),
    .A3(_11333_),
    .ZN(_11409_));
 NOR2_X1 _35314_ (.A1(_11328_),
    .A2(_11293_),
    .ZN(_11410_));
 NAND4_X1 _35315_ (.A1(_20636_),
    .A2(_11408_),
    .A3(_11409_),
    .A4(_11410_),
    .ZN(_11411_));
 OAI21_X1 _35316_ (.A(_11319_),
    .B1(_11295_),
    .B2(_11294_),
    .ZN(_11412_));
 NAND3_X1 _35317_ (.A1(_11215_),
    .A2(_11219_),
    .A3(_11261_),
    .ZN(_11413_));
 OAI221_X2 _35318_ (.A(_11412_),
    .B1(_11413_),
    .B2(_11290_),
    .C1(_11258_),
    .C2(_11264_),
    .ZN(_11414_));
 NAND4_X1 _35319_ (.A1(_11338_),
    .A2(_11368_),
    .A3(_20636_),
    .A4(_11414_),
    .ZN(_11415_));
 NAND2_X1 _35320_ (.A1(_11194_),
    .A2(_11299_),
    .ZN(_11416_));
 AOI21_X1 _35321_ (.A(_11416_),
    .B1(_11325_),
    .B2(_11331_),
    .ZN(_11417_));
 OAI21_X1 _35322_ (.A(_11315_),
    .B1(_11302_),
    .B2(_11304_),
    .ZN(_11418_));
 AOI221_X1 _35323_ (.A(_11417_),
    .B1(_11418_),
    .B2(_11194_),
    .C1(_20614_),
    .C2(_11301_),
    .ZN(_11419_));
 NAND3_X1 _35324_ (.A1(_11411_),
    .A2(_11415_),
    .A3(_11419_),
    .ZN(_11420_));
 NAND2_X1 _35325_ (.A1(_11368_),
    .A2(_11301_),
    .ZN(_11421_));
 AOI21_X1 _35326_ (.A(_11266_),
    .B1(_11361_),
    .B2(_11371_),
    .ZN(_11422_));
 NAND3_X1 _35327_ (.A1(_11215_),
    .A2(_11219_),
    .A3(_11253_),
    .ZN(_11423_));
 OAI21_X1 _35328_ (.A(_11330_),
    .B1(_11331_),
    .B2(_11423_),
    .ZN(_11424_));
 AOI21_X2 _35329_ (.A(_11235_),
    .B1(_11245_),
    .B2(_11371_),
    .ZN(_11425_));
 NAND2_X1 _35330_ (.A1(_11242_),
    .A2(_11245_),
    .ZN(_11426_));
 OAI21_X1 _35331_ (.A(_11338_),
    .B1(_11375_),
    .B2(_11426_),
    .ZN(_11427_));
 OAI22_X2 _35332_ (.A1(_11422_),
    .A2(_11424_),
    .B1(_11425_),
    .B2(_11427_),
    .ZN(_11428_));
 NAND2_X1 _35333_ (.A1(_11338_),
    .A2(_11225_),
    .ZN(_11429_));
 NAND3_X1 _35334_ (.A1(_11215_),
    .A2(_11219_),
    .A3(_11232_),
    .ZN(_11430_));
 NOR3_X1 _35335_ (.A1(_11294_),
    .A2(_11295_),
    .A3(_11225_),
    .ZN(_11431_));
 OAI21_X2 _35336_ (.A(_11430_),
    .B1(_11431_),
    .B2(_11228_),
    .ZN(_11432_));
 OAI221_X2 _35337_ (.A(_11368_),
    .B1(_11375_),
    .B2(_11429_),
    .C1(_11432_),
    .C2(_11338_),
    .ZN(_11433_));
 OAI221_X2 _35338_ (.A(_20641_),
    .B1(_11421_),
    .B2(_11428_),
    .C1(_11433_),
    .C2(_11301_),
    .ZN(_11434_));
 NAND3_X1 _35339_ (.A1(_11371_),
    .A2(_11420_),
    .A3(_11434_),
    .ZN(_11435_));
 AND2_X1 _35340_ (.A1(_11367_),
    .A2(_11368_),
    .ZN(_11436_));
 NAND3_X1 _35341_ (.A1(_11368_),
    .A2(_11420_),
    .A3(_11434_),
    .ZN(_11437_));
 NOR2_X1 _35342_ (.A1(_11367_),
    .A2(_11375_),
    .ZN(_11438_));
 AOI22_X2 _35343_ (.A1(_11435_),
    .A2(_11436_),
    .B1(_11437_),
    .B2(_11438_),
    .ZN(_11439_));
 OAI21_X1 _35344_ (.A(_11330_),
    .B1(_11375_),
    .B2(_11426_),
    .ZN(_11440_));
 OAI22_X2 _35345_ (.A1(_11330_),
    .A2(_11432_),
    .B1(_11440_),
    .B2(_11425_),
    .ZN(_11441_));
 MUX2_X1 _35346_ (.A(_11228_),
    .B(_11225_),
    .S(_11308_),
    .Z(_11442_));
 OAI22_X2 _35347_ (.A1(_11327_),
    .A2(_11441_),
    .B1(_11442_),
    .B2(_11314_),
    .ZN(_11443_));
 AOI21_X1 _35348_ (.A(_11305_),
    .B1(_11325_),
    .B2(_11299_),
    .ZN(_11444_));
 NOR2_X1 _35349_ (.A1(_20611_),
    .A2(_11444_),
    .ZN(_11445_));
 MUX2_X1 _35350_ (.A(_11300_),
    .B(_11445_),
    .S(_11291_),
    .Z(_11446_));
 AOI22_X2 _35351_ (.A1(_20613_),
    .A2(_11335_),
    .B1(_11334_),
    .B2(_11314_),
    .ZN(_11447_));
 NOR2_X1 _35352_ (.A1(_11418_),
    .A2(_11447_),
    .ZN(_11448_));
 MUX2_X1 _35353_ (.A(_11266_),
    .B(_11258_),
    .S(_11329_),
    .Z(_11449_));
 NAND2_X1 _35354_ (.A1(_11194_),
    .A2(_11449_),
    .ZN(_11450_));
 AND2_X1 _35355_ (.A1(_11331_),
    .A2(_11450_),
    .ZN(_11451_));
 AOI21_X1 _35356_ (.A(_11331_),
    .B1(_11387_),
    .B2(_11371_),
    .ZN(_11452_));
 OAI222_X2 _35357_ (.A1(_11194_),
    .A2(_11378_),
    .B1(_11451_),
    .B2(_11452_),
    .C1(_11450_),
    .C2(_11371_),
    .ZN(_11453_));
 INV_X1 _35358_ (.A(_11453_),
    .ZN(_11454_));
 AND2_X1 _35359_ (.A1(_20641_),
    .A2(_11405_),
    .ZN(_11455_));
 AOI221_X2 _35360_ (.A(_11443_),
    .B1(_11446_),
    .B2(_11448_),
    .C1(_11454_),
    .C2(_11455_),
    .ZN(_11456_));
 NAND2_X1 _35361_ (.A1(_11329_),
    .A2(_11253_),
    .ZN(_11457_));
 NAND2_X1 _35362_ (.A1(_11328_),
    .A2(_11242_),
    .ZN(_11458_));
 AOI22_X2 _35363_ (.A1(_11371_),
    .A2(_11361_),
    .B1(_11457_),
    .B2(_11458_),
    .ZN(_11459_));
 NOR4_X2 _35364_ (.A1(_11338_),
    .A2(_11220_),
    .A3(_11258_),
    .A4(_11331_),
    .ZN(_11460_));
 NOR4_X2 _35365_ (.A1(_11329_),
    .A2(_11220_),
    .A3(_11266_),
    .A4(_11331_),
    .ZN(_11461_));
 NOR3_X2 _35366_ (.A1(_11459_),
    .A2(_11460_),
    .A3(_11461_),
    .ZN(_11462_));
 INV_X1 _35367_ (.A(_11291_),
    .ZN(_11463_));
 NOR2_X1 _35368_ (.A1(_11463_),
    .A2(_11315_),
    .ZN(_11464_));
 NAND2_X1 _35369_ (.A1(_11463_),
    .A2(_11299_),
    .ZN(_11465_));
 AOI21_X2 _35370_ (.A(_11465_),
    .B1(_11325_),
    .B2(_11290_),
    .ZN(_11466_));
 OAI21_X4 _35371_ (.A(_11314_),
    .B1(_11464_),
    .B2(_11466_),
    .ZN(_11467_));
 NOR2_X1 _35372_ (.A1(_11462_),
    .A2(_11467_),
    .ZN(_11468_));
 MUX2_X1 _35373_ (.A(_11296_),
    .B(_11375_),
    .S(_11367_),
    .Z(_11469_));
 AOI21_X2 _35374_ (.A(_11468_),
    .B1(_11469_),
    .B2(_11306_),
    .ZN(_11470_));
 NAND2_X1 _35375_ (.A1(_11330_),
    .A2(_11401_),
    .ZN(_11471_));
 NAND2_X1 _35376_ (.A1(_11338_),
    .A2(_11296_),
    .ZN(_11472_));
 OAI21_X1 _35377_ (.A(_11471_),
    .B1(_11472_),
    .B2(_11373_),
    .ZN(_11473_));
 AND2_X1 _35378_ (.A1(_11244_),
    .A2(_11374_),
    .ZN(_11474_));
 OR2_X1 _35379_ (.A1(_11220_),
    .A2(_11335_),
    .ZN(_11475_));
 NAND2_X1 _35380_ (.A1(_11296_),
    .A2(_11311_),
    .ZN(_11476_));
 MUX2_X1 _35381_ (.A(_11261_),
    .B(_11476_),
    .S(_11214_),
    .Z(_11477_));
 MUX2_X1 _35382_ (.A(_11261_),
    .B(_11476_),
    .S(_11213_),
    .Z(_11478_));
 NOR2_X1 _35383_ (.A1(_11218_),
    .A2(_11130_),
    .ZN(_11479_));
 MUX2_X1 _35384_ (.A(_11477_),
    .B(_11478_),
    .S(_11479_),
    .Z(_11480_));
 OAI221_X2 _35385_ (.A(_11194_),
    .B1(_11474_),
    .B2(_11475_),
    .C1(_11480_),
    .C2(_11330_),
    .ZN(_11481_));
 NAND3_X1 _35386_ (.A1(_11338_),
    .A2(_11385_),
    .A3(_11331_),
    .ZN(_11482_));
 OAI21_X2 _35387_ (.A(_11482_),
    .B1(_11339_),
    .B2(_11338_),
    .ZN(_11483_));
 NOR3_X1 _35388_ (.A1(_20641_),
    .A2(_11481_),
    .A3(_11483_),
    .ZN(_11484_));
 OAI21_X2 _35389_ (.A(_11392_),
    .B1(_11473_),
    .B2(_11484_),
    .ZN(_11485_));
 AOI21_X2 _35390_ (.A(_11456_),
    .B1(_11470_),
    .B2(_11485_),
    .ZN(_11486_));
 NAND2_X1 _35391_ (.A1(_11308_),
    .A2(_11228_),
    .ZN(_11487_));
 OAI221_X2 _35392_ (.A(_11487_),
    .B1(_11375_),
    .B2(_11293_),
    .C1(_11367_),
    .C2(_11232_),
    .ZN(_11488_));
 OAI21_X2 _35393_ (.A(_11488_),
    .B1(_11467_),
    .B2(_11390_),
    .ZN(_11489_));
 AOI21_X4 _35394_ (.A(_11489_),
    .B1(_11392_),
    .B2(_11404_),
    .ZN(_11490_));
 INV_X1 _35395_ (.A(_11490_),
    .ZN(_11491_));
 MUX2_X1 _35396_ (.A(_11235_),
    .B(_11400_),
    .S(_11307_),
    .Z(_11492_));
 NOR2_X1 _35397_ (.A1(_11314_),
    .A2(_11492_),
    .ZN(_11493_));
 NAND2_X1 _35398_ (.A1(_20613_),
    .A2(_11380_),
    .ZN(_11494_));
 OR3_X1 _35399_ (.A1(_11338_),
    .A2(_20613_),
    .A3(_11333_),
    .ZN(_11495_));
 MUX2_X1 _35400_ (.A(_11258_),
    .B(_11385_),
    .S(_20611_),
    .Z(_11496_));
 OAI211_X2 _35401_ (.A(_11494_),
    .B(_11495_),
    .C1(_11496_),
    .C2(_11330_),
    .ZN(_11497_));
 INV_X1 _35402_ (.A(_20614_),
    .ZN(_11498_));
 OAI21_X1 _35403_ (.A(_11428_),
    .B1(_20641_),
    .B2(_11498_),
    .ZN(_11499_));
 AOI221_X2 _35404_ (.A(_11493_),
    .B1(_11497_),
    .B2(_11455_),
    .C1(_11392_),
    .C2(_11499_),
    .ZN(_11500_));
 NOR2_X1 _35405_ (.A1(_11307_),
    .A2(_11266_),
    .ZN(_11501_));
 AOI21_X1 _35406_ (.A(_11501_),
    .B1(_11242_),
    .B2(_11308_),
    .ZN(_11502_));
 OAI222_X2 _35407_ (.A1(_11467_),
    .A2(_11447_),
    .B1(_11453_),
    .B2(_11327_),
    .C1(_11314_),
    .C2(_11502_),
    .ZN(_11503_));
 INV_X1 _35408_ (.A(_11503_),
    .ZN(_11504_));
 MUX2_X1 _35409_ (.A(_11385_),
    .B(_11258_),
    .S(_11307_),
    .Z(_11505_));
 OAI33_X1 _35410_ (.A1(_11327_),
    .A2(_11481_),
    .A3(_11483_),
    .B1(_11505_),
    .B2(_11302_),
    .B3(_11304_),
    .ZN(_20618_));
 NAND3_X2 _35411_ (.A1(_11337_),
    .A2(_11342_),
    .A3(_20618_),
    .ZN(_11506_));
 NOR2_X1 _35412_ (.A1(_11307_),
    .A2(_11258_),
    .ZN(_11507_));
 AOI221_X2 _35413_ (.A(_11507_),
    .B1(_11370_),
    .B2(_11194_),
    .C1(_11307_),
    .C2(_11253_),
    .ZN(_11508_));
 OAI21_X1 _35414_ (.A(_11290_),
    .B1(_11305_),
    .B2(_11325_),
    .ZN(_11509_));
 AOI211_X2 _35415_ (.A(_11297_),
    .B(_11305_),
    .C1(_11509_),
    .C2(_11299_),
    .ZN(_11510_));
 OAI221_X1 _35416_ (.A(_11291_),
    .B1(_11297_),
    .B2(_11298_),
    .C1(_11302_),
    .C2(_11304_),
    .ZN(_11511_));
 OR3_X1 _35417_ (.A1(_11291_),
    .A2(_11302_),
    .A3(_11304_),
    .ZN(_11512_));
 AND4_X1 _35418_ (.A1(_11328_),
    .A2(_11465_),
    .A3(_11511_),
    .A4(_11512_),
    .ZN(_11513_));
 AOI221_X1 _35419_ (.A(_11305_),
    .B1(_11414_),
    .B2(_11513_),
    .C1(_11301_),
    .C2(_20614_),
    .ZN(_11514_));
 AOI211_X4 _35420_ (.A(_11508_),
    .B(_11510_),
    .C1(_11514_),
    .C2(_11411_),
    .ZN(_11515_));
 MUX2_X1 _35421_ (.A(_11253_),
    .B(_11250_),
    .S(_11307_),
    .Z(_11516_));
 NAND2_X1 _35422_ (.A1(_11305_),
    .A2(_11516_),
    .ZN(_11517_));
 OAI221_X1 _35423_ (.A(_11517_),
    .B1(_11467_),
    .B2(_11340_),
    .C1(_11327_),
    .C2(_11390_),
    .ZN(_11518_));
 NOR3_X2 _35424_ (.A1(_11481_),
    .A2(_11483_),
    .A3(_11467_),
    .ZN(_11519_));
 NAND2_X1 _35425_ (.A1(_11308_),
    .A2(_11235_),
    .ZN(_11520_));
 OAI221_X2 _35426_ (.A(_11520_),
    .B1(_11375_),
    .B2(_11293_),
    .C1(_11308_),
    .C2(_11242_),
    .ZN(_11521_));
 OAI21_X2 _35427_ (.A(_11521_),
    .B1(_11462_),
    .B2(_11327_),
    .ZN(_11522_));
 OAI211_X4 _35428_ (.A(_11515_),
    .B(_11518_),
    .C1(_11519_),
    .C2(_11522_),
    .ZN(_11523_));
 NOR4_X1 _35429_ (.A1(_11500_),
    .A2(_11504_),
    .A3(_11506_),
    .A4(_11523_),
    .ZN(_11524_));
 NAND4_X2 _35430_ (.A1(_11439_),
    .A2(_11486_),
    .A3(_11491_),
    .A4(_11524_),
    .ZN(_11525_));
 XNOR2_X1 _35431_ (.A(_11407_),
    .B(_11525_),
    .ZN(_11526_));
 MUX2_X1 _35432_ (.A(_11348_),
    .B(_11366_),
    .S(_11526_),
    .Z(_11527_));
 NAND2_X2 _35433_ (.A1(_10973_),
    .A2(_11345_),
    .ZN(_11528_));
 OAI21_X1 _35434_ (.A(_11347_),
    .B1(_11527_),
    .B2(_11528_),
    .ZN(_00016_));
 CLKBUF_X3 _35435_ (.A(_10973_),
    .Z(_11529_));
 NAND2_X4 _35436_ (.A1(_10973_),
    .A2(_10976_),
    .ZN(_11530_));
 OAI22_X1 _35437_ (.A1(\g_reduce0[10].adder.b[1] ),
    .A2(_11529_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[1] ),
    .ZN(_11531_));
 XOR2_X1 _35438_ (.A(_20620_),
    .B(_11515_),
    .Z(_11532_));
 NOR2_X1 _35439_ (.A1(_11528_),
    .A2(_11532_),
    .ZN(_11533_));
 NOR2_X1 _35440_ (.A1(_20621_),
    .A2(_11528_),
    .ZN(_11534_));
 MUX2_X1 _35441_ (.A(_11533_),
    .B(_11534_),
    .S(_11526_),
    .Z(_11535_));
 NOR2_X1 _35442_ (.A1(_11531_),
    .A2(_11535_),
    .ZN(_00023_));
 OAI22_X2 _35443_ (.A1(\g_reduce0[10].adder.b[2] ),
    .A2(_10973_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[2] ),
    .ZN(_11536_));
 AND3_X1 _35444_ (.A1(_20619_),
    .A2(_11515_),
    .A3(_20618_),
    .ZN(_11537_));
 XNOR2_X1 _35445_ (.A(_11518_),
    .B(_11537_),
    .ZN(_11538_));
 NOR2_X1 _35446_ (.A1(_11343_),
    .A2(_10976_),
    .ZN(_11539_));
 AOI21_X1 _35447_ (.A(_11536_),
    .B1(_11538_),
    .B2(_11539_),
    .ZN(_11540_));
 NOR2_X1 _35448_ (.A1(_11533_),
    .A2(_11536_),
    .ZN(_11541_));
 MUX2_X1 _35449_ (.A(_11540_),
    .B(_11541_),
    .S(_11526_),
    .Z(_00024_));
 AOI22_X1 _35450_ (.A1(\g_reduce0[10].adder.b[3] ),
    .A2(_11343_),
    .B1(_11346_),
    .B2(\g_reduce0[10].adder.a[3] ),
    .ZN(_11542_));
 AND2_X1 _35451_ (.A1(_11515_),
    .A2(_11518_),
    .ZN(_11543_));
 NAND2_X1 _35452_ (.A1(_20620_),
    .A2(_11543_),
    .ZN(_11544_));
 XNOR2_X1 _35453_ (.A(_11504_),
    .B(_11544_),
    .ZN(_11545_));
 MUX2_X1 _35454_ (.A(_11545_),
    .B(_11538_),
    .S(_11526_),
    .Z(_11546_));
 OAI21_X1 _35455_ (.A(_11542_),
    .B1(_11546_),
    .B2(_11528_),
    .ZN(_00025_));
 OAI22_X1 _35456_ (.A1(\g_reduce0[10].adder.b[4] ),
    .A2(_11529_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[4] ),
    .ZN(_11547_));
 NOR2_X1 _35457_ (.A1(_11519_),
    .A2(_11522_),
    .ZN(_11548_));
 NAND2_X1 _35458_ (.A1(_11503_),
    .A2(_11543_),
    .ZN(_11549_));
 NOR2_X1 _35459_ (.A1(_11549_),
    .A2(_11506_),
    .ZN(_11550_));
 XOR2_X1 _35460_ (.A(_11548_),
    .B(_11550_),
    .Z(_11551_));
 MUX2_X1 _35461_ (.A(_11551_),
    .B(_11545_),
    .S(_11526_),
    .Z(_11552_));
 AOI21_X1 _35462_ (.A(_11547_),
    .B1(_11552_),
    .B2(_11539_),
    .ZN(_00026_));
 AOI22_X1 _35463_ (.A1(\g_reduce0[10].adder.b[5] ),
    .A2(_11343_),
    .B1(_11346_),
    .B2(\g_reduce0[10].adder.a[5] ),
    .ZN(_11553_));
 NAND2_X1 _35464_ (.A1(_11455_),
    .A2(_11497_),
    .ZN(_11554_));
 AOI21_X1 _35465_ (.A(_11493_),
    .B1(_11499_),
    .B2(_11392_),
    .ZN(_11555_));
 NAND2_X1 _35466_ (.A1(_11554_),
    .A2(_11555_),
    .ZN(_11556_));
 NAND2_X2 _35467_ (.A1(_20620_),
    .A2(_11503_),
    .ZN(_11557_));
 NOR2_X1 _35468_ (.A1(_11523_),
    .A2(_11557_),
    .ZN(_11558_));
 XNOR2_X1 _35469_ (.A(_11556_),
    .B(_11558_),
    .ZN(_11559_));
 MUX2_X1 _35470_ (.A(_11559_),
    .B(_11551_),
    .S(_11526_),
    .Z(_11560_));
 OAI21_X1 _35471_ (.A(_11553_),
    .B1(_11560_),
    .B2(_11528_),
    .ZN(_00027_));
 OAI21_X1 _35472_ (.A(_11500_),
    .B1(_11523_),
    .B2(_11557_),
    .ZN(_11561_));
 OAI22_X2 _35473_ (.A1(\g_reduce0[10].adder.b[6] ),
    .A2(_10973_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[6] ),
    .ZN(_11562_));
 AOI21_X1 _35474_ (.A(_11562_),
    .B1(_11558_),
    .B2(_11556_),
    .ZN(_11563_));
 NAND3_X1 _35475_ (.A1(_11526_),
    .A2(_11561_),
    .A3(_11563_),
    .ZN(_11564_));
 XNOR2_X1 _35476_ (.A(_11491_),
    .B(_11524_),
    .ZN(_11565_));
 NOR2_X1 _35477_ (.A1(_11407_),
    .A2(_11565_),
    .ZN(_11566_));
 NOR2_X1 _35478_ (.A1(_11528_),
    .A2(_11566_),
    .ZN(_11567_));
 OAI21_X1 _35479_ (.A(_11564_),
    .B1(_11567_),
    .B2(_11562_),
    .ZN(_00028_));
 NAND3_X2 _35480_ (.A1(_11369_),
    .A2(_11393_),
    .A3(_11406_),
    .ZN(_11568_));
 OAI21_X1 _35481_ (.A(_11539_),
    .B1(_11568_),
    .B2(_11565_),
    .ZN(_11569_));
 OAI221_X1 _35482_ (.A(_11569_),
    .B1(_11529_),
    .B2(\g_reduce0[10].adder.b[7] ),
    .C1(\g_reduce0[10].adder.a[7] ),
    .C2(_11530_),
    .ZN(_11570_));
 NOR4_X4 _35483_ (.A1(_11500_),
    .A2(_11490_),
    .A3(_11523_),
    .A4(_11557_),
    .ZN(_11571_));
 XNOR2_X1 _35484_ (.A(_11456_),
    .B(_11571_),
    .ZN(_11572_));
 OAI221_X1 _35485_ (.A(_11572_),
    .B1(_11529_),
    .B2(\g_reduce0[10].adder.b[7] ),
    .C1(\g_reduce0[10].adder.a[7] ),
    .C2(_11530_),
    .ZN(_11573_));
 OAI21_X1 _35486_ (.A(_11570_),
    .B1(_11573_),
    .B2(_11526_),
    .ZN(_00029_));
 OAI22_X1 _35487_ (.A1(\g_reduce0[10].adder.b[8] ),
    .A2(_11529_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[8] ),
    .ZN(_11574_));
 AND3_X1 _35488_ (.A1(_11486_),
    .A2(_11491_),
    .A3(_11524_),
    .ZN(_11575_));
 NAND2_X1 _35489_ (.A1(_11485_),
    .A2(_11470_),
    .ZN(_11576_));
 NOR2_X1 _35490_ (.A1(_11456_),
    .A2(_11490_),
    .ZN(_11577_));
 AOI21_X1 _35491_ (.A(_11576_),
    .B1(_11524_),
    .B2(_11577_),
    .ZN(_11578_));
 NOR3_X1 _35492_ (.A1(_11407_),
    .A2(_11575_),
    .A3(_11578_),
    .ZN(_11579_));
 NOR2_X1 _35493_ (.A1(_11528_),
    .A2(_11579_),
    .ZN(_11580_));
 NAND2_X1 _35494_ (.A1(_11526_),
    .A2(_11572_),
    .ZN(_11581_));
 AOI21_X1 _35495_ (.A(_11574_),
    .B1(_11580_),
    .B2(_11581_),
    .ZN(_00030_));
 OAI22_X2 _35496_ (.A1(\g_reduce0[10].adder.b[9] ),
    .A2(_10973_),
    .B1(_11530_),
    .B2(\g_reduce0[10].adder.a[9] ),
    .ZN(_11582_));
 AND3_X1 _35497_ (.A1(_11371_),
    .A2(_11420_),
    .A3(_11434_),
    .ZN(_11583_));
 NAND2_X1 _35498_ (.A1(_11367_),
    .A2(_11368_),
    .ZN(_11584_));
 AND3_X1 _35499_ (.A1(_11368_),
    .A2(_11420_),
    .A3(_11434_),
    .ZN(_11585_));
 OR2_X1 _35500_ (.A1(_11367_),
    .A2(_11375_),
    .ZN(_11586_));
 OAI22_X4 _35501_ (.A1(_11583_),
    .A2(_11584_),
    .B1(_11585_),
    .B2(_11586_),
    .ZN(_11587_));
 NOR2_X1 _35502_ (.A1(_11587_),
    .A2(_11571_),
    .ZN(_11588_));
 AOI21_X1 _35503_ (.A(_11407_),
    .B1(_11491_),
    .B2(_11524_),
    .ZN(_11589_));
 NOR2_X1 _35504_ (.A1(_11568_),
    .A2(_11587_),
    .ZN(_11590_));
 NOR3_X1 _35505_ (.A1(_11407_),
    .A2(_11439_),
    .A3(_11456_),
    .ZN(_11591_));
 MUX2_X1 _35506_ (.A(_11590_),
    .B(_11591_),
    .S(_11571_),
    .Z(_11592_));
 AOI221_X1 _35507_ (.A(_11528_),
    .B1(_11588_),
    .B2(_11589_),
    .C1(_11592_),
    .C2(_11576_),
    .ZN(_11593_));
 OAI21_X1 _35508_ (.A(_11568_),
    .B1(_11587_),
    .B2(_11486_),
    .ZN(_11594_));
 NAND3_X1 _35509_ (.A1(_11407_),
    .A2(_11485_),
    .A3(_11470_),
    .ZN(_11595_));
 AND2_X1 _35510_ (.A1(_11524_),
    .A2(_11577_),
    .ZN(_11596_));
 OAI21_X1 _35511_ (.A(_11594_),
    .B1(_11595_),
    .B2(_11596_),
    .ZN(_11597_));
 OR2_X1 _35512_ (.A1(_11575_),
    .A2(_11582_),
    .ZN(_11598_));
 OAI22_X1 _35513_ (.A1(_11582_),
    .A2(_11593_),
    .B1(_11597_),
    .B2(_11598_),
    .ZN(_00031_));
 INV_X1 _35514_ (.A(_20628_),
    .ZN(_20622_));
 MUX2_X1 _35515_ (.A(\g_reduce0[10].adder.a[10] ),
    .B(_20627_),
    .S(_11345_),
    .Z(_11599_));
 MUX2_X1 _35516_ (.A(\g_reduce0[10].adder.b[10] ),
    .B(_11599_),
    .S(_11529_),
    .Z(_00017_));
 MUX2_X1 _35517_ (.A(\g_reduce0[10].adder.a[11] ),
    .B(_20635_),
    .S(_11345_),
    .Z(_11600_));
 MUX2_X1 _35518_ (.A(\g_reduce0[10].adder.b[11] ),
    .B(_11600_),
    .S(_11529_),
    .Z(_00018_));
 XOR2_X1 _35519_ (.A(_14519_),
    .B(_20639_),
    .Z(_11601_));
 MUX2_X1 _35520_ (.A(_20503_),
    .B(_00472_),
    .S(_11023_),
    .Z(_11602_));
 NAND2_X1 _35521_ (.A1(_11308_),
    .A2(_20629_),
    .ZN(_11603_));
 XOR2_X1 _35522_ (.A(_11602_),
    .B(_11603_),
    .Z(_11604_));
 MUX2_X1 _35523_ (.A(_11601_),
    .B(_11604_),
    .S(_11306_),
    .Z(_11605_));
 XOR2_X1 _35524_ (.A(_20634_),
    .B(_11605_),
    .Z(_11606_));
 MUX2_X1 _35525_ (.A(\g_reduce0[10].adder.a[12] ),
    .B(_11606_),
    .S(_11345_),
    .Z(_11607_));
 MUX2_X1 _35526_ (.A(\g_reduce0[10].adder.b[12] ),
    .B(_11607_),
    .S(_11529_),
    .Z(_00019_));
 INV_X1 _35527_ (.A(_14521_),
    .ZN(_14518_));
 INV_X1 _35528_ (.A(_20631_),
    .ZN(_11608_));
 INV_X1 _35529_ (.A(_20632_),
    .ZN(_11609_));
 OAI21_X1 _35530_ (.A(_11608_),
    .B1(_11609_),
    .B2(_14521_),
    .ZN(_11610_));
 AOI21_X1 _35531_ (.A(_20638_),
    .B1(_11610_),
    .B2(_20639_),
    .ZN(_11611_));
 XNOR2_X1 _35532_ (.A(_20643_),
    .B(_11611_),
    .ZN(_11612_));
 MUX2_X1 _35533_ (.A(_20500_),
    .B(_00475_),
    .S(_11023_),
    .Z(_11613_));
 INV_X1 _35534_ (.A(_11602_),
    .ZN(_20637_));
 MUX2_X1 _35535_ (.A(_20506_),
    .B(_00467_),
    .S(_11023_),
    .Z(_11614_));
 INV_X2 _35536_ (.A(_11614_),
    .ZN(_14516_));
 AND4_X1 _35537_ (.A1(_11308_),
    .A2(_20628_),
    .A3(_20637_),
    .A4(_14516_),
    .ZN(_11615_));
 XNOR2_X1 _35538_ (.A(_11613_),
    .B(_11615_),
    .ZN(_11616_));
 MUX2_X1 _35539_ (.A(_11612_),
    .B(_11616_),
    .S(_11306_),
    .Z(_11617_));
 NAND2_X1 _35540_ (.A1(_11367_),
    .A2(_20630_),
    .ZN(_11618_));
 OAI21_X1 _35541_ (.A(_11618_),
    .B1(_11614_),
    .B2(_11367_),
    .ZN(_11619_));
 MUX2_X1 _35542_ (.A(_14520_),
    .B(_11619_),
    .S(_11306_),
    .Z(_20633_));
 NAND3_X1 _35543_ (.A1(_20626_),
    .A2(_11605_),
    .A3(_20633_),
    .ZN(_11620_));
 XNOR2_X1 _35544_ (.A(_11617_),
    .B(_11620_),
    .ZN(_11621_));
 MUX2_X1 _35545_ (.A(\g_reduce0[10].adder.a[13] ),
    .B(_11621_),
    .S(_11345_),
    .Z(_11622_));
 MUX2_X1 _35546_ (.A(\g_reduce0[10].adder.b[13] ),
    .B(_11622_),
    .S(_11529_),
    .Z(_00020_));
 OR2_X1 _35547_ (.A1(_10974_),
    .A2(_11012_),
    .ZN(_11623_));
 NAND2_X1 _35548_ (.A1(\g_reduce0[10].adder.a[14] ),
    .A2(_11623_),
    .ZN(_11624_));
 NOR4_X1 _35549_ (.A1(_11314_),
    .A2(_11602_),
    .A3(_11603_),
    .A4(_11613_),
    .ZN(_11625_));
 AOI21_X1 _35550_ (.A(_20638_),
    .B1(_20639_),
    .B2(_14519_),
    .ZN(_11626_));
 INV_X1 _35551_ (.A(_11626_),
    .ZN(_11627_));
 AOI21_X1 _35552_ (.A(_20642_),
    .B1(_11627_),
    .B2(_20643_),
    .ZN(_11628_));
 AOI21_X2 _35553_ (.A(_11625_),
    .B1(_11628_),
    .B2(_11314_),
    .ZN(_11629_));
 NAND3_X1 _35554_ (.A1(_20634_),
    .A2(_11605_),
    .A3(_11617_),
    .ZN(_11630_));
 XNOR2_X2 _35555_ (.A(_11629_),
    .B(_11630_),
    .ZN(_11631_));
 MUX2_X1 _35556_ (.A(_11624_),
    .B(_11623_),
    .S(_11631_),
    .Z(_11632_));
 OAI22_X1 _35557_ (.A1(_10974_),
    .A2(_11529_),
    .B1(_10976_),
    .B2(_11632_),
    .ZN(_11633_));
 NOR2_X1 _35558_ (.A1(\g_reduce0[10].adder.a[14] ),
    .A2(_11343_),
    .ZN(_11634_));
 AOI21_X1 _35559_ (.A(_10976_),
    .B1(_11012_),
    .B2(_11631_),
    .ZN(_11635_));
 NAND2_X1 _35560_ (.A1(_10974_),
    .A2(_11060_),
    .ZN(_11636_));
 OAI21_X1 _35561_ (.A(_11635_),
    .B1(_11636_),
    .B2(_11631_),
    .ZN(_11637_));
 AOI21_X1 _35562_ (.A(_11633_),
    .B1(_11634_),
    .B2(_11637_),
    .ZN(_00021_));
 BUF_X1 _35563_ (.A(b[15]),
    .Z(_11638_));
 XOR2_X1 _35564_ (.A(_11638_),
    .B(net60),
    .Z(_00207_));
 BUF_X1 _35565_ (.A(b[31]),
    .Z(_11639_));
 XOR2_X1 _35566_ (.A(_11639_),
    .B(net162),
    .Z(_00223_));
 BUF_X1 _35567_ (.A(b[47]),
    .Z(_11640_));
 XOR2_X1 _35568_ (.A(_11640_),
    .B(net178),
    .Z(_00239_));
 BUF_X1 _35569_ (.A(b[63]),
    .Z(_11641_));
 XOR2_X1 _35570_ (.A(_11641_),
    .B(net194),
    .Z(_00255_));
 XOR2_X1 _35571_ (.A(_11638_),
    .B(net210),
    .Z(_00271_));
 XOR2_X1 _35572_ (.A(_11639_),
    .B(net227),
    .Z(_00287_));
 XOR2_X1 _35573_ (.A(_11640_),
    .B(net12),
    .Z(_00303_));
 XOR2_X1 _35574_ (.A(_11641_),
    .B(net27),
    .Z(_00319_));
 XOR2_X1 _35575_ (.A(_11638_),
    .B(net43),
    .Z(_00335_));
 XOR2_X1 _35576_ (.A(_11639_),
    .B(net59),
    .Z(_00351_));
 XOR2_X1 _35577_ (.A(_11640_),
    .B(net75),
    .Z(_00367_));
 XOR2_X1 _35578_ (.A(_11641_),
    .B(net91),
    .Z(_00383_));
 XOR2_X1 _35579_ (.A(_11638_),
    .B(net107),
    .Z(_00399_));
 XOR2_X1 _35580_ (.A(_11639_),
    .B(net124),
    .Z(_00415_));
 XOR2_X1 _35581_ (.A(_11640_),
    .B(net140),
    .Z(_00431_));
 XOR2_X1 _35582_ (.A(_11641_),
    .B(net155),
    .Z(_00447_));
 BUF_X1 _35583_ (.A(net28),
    .Z(_11642_));
 BUF_X1 _35584_ (.A(b[9]),
    .Z(_11643_));
 AND2_X1 _35585_ (.A1(_11642_),
    .A2(_11643_),
    .ZN(_20644_));
 BUF_X2 _35586_ (.A(net29),
    .Z(_11644_));
 BUF_X1 _35587_ (.A(net275),
    .Z(_11645_));
 AND2_X1 _35588_ (.A1(_11644_),
    .A2(_11645_),
    .ZN(_20645_));
 BUF_X2 _35589_ (.A(net33),
    .Z(_11646_));
 BUF_X1 _35590_ (.A(net270),
    .Z(_11647_));
 BUF_X1 _35591_ (.A(_11647_),
    .Z(_11648_));
 AND2_X1 _35592_ (.A1(_11646_),
    .A2(_11648_),
    .ZN(_14529_));
 BUF_X2 _35593_ (.A(net31),
    .Z(_11649_));
 BUF_X1 _35594_ (.A(net274),
    .Z(_11650_));
 CLKBUF_X3 _35595_ (.A(_11650_),
    .Z(_11651_));
 AND2_X1 _35596_ (.A1(_11649_),
    .A2(_11651_),
    .ZN(_14528_));
 BUF_X2 _35597_ (.A(net32),
    .Z(_11652_));
 CLKBUF_X3 _35598_ (.A(b[6]),
    .Z(_11653_));
 BUF_X2 _35599_ (.A(_11653_),
    .Z(_11654_));
 AND2_X1 _35600_ (.A1(_11652_),
    .A2(_11654_),
    .ZN(_14527_));
 BUF_X2 _35601_ (.A(a[135]),
    .Z(_11655_));
 BUF_X1 _35602_ (.A(net248),
    .Z(_11656_));
 BUF_X1 _35603_ (.A(_11656_),
    .Z(_11657_));
 AND2_X1 _35604_ (.A1(_11655_),
    .A2(_11657_),
    .ZN(_14532_));
 BUF_X2 _35605_ (.A(net34),
    .Z(_11658_));
 BUF_X1 _35606_ (.A(net262),
    .Z(_11659_));
 BUF_X2 _35607_ (.A(_11659_),
    .Z(_11660_));
 AND2_X1 _35608_ (.A1(_11658_),
    .A2(_11660_),
    .ZN(_14533_));
 BUF_X2 _35609_ (.A(net35),
    .Z(_11661_));
 CLKBUF_X3 _35610_ (.A(b[3]),
    .Z(_11662_));
 BUF_X2 _35611_ (.A(_11662_),
    .Z(_11663_));
 AND2_X1 _35612_ (.A1(_11661_),
    .A2(_11663_),
    .ZN(_14534_));
 BUF_X1 _35613_ (.A(_11656_),
    .Z(_11664_));
 AND2_X1 _35614_ (.A1(_11664_),
    .A2(_11661_),
    .ZN(_20650_));
 BUF_X4 _35615_ (.A(b[1]),
    .Z(_11665_));
 INV_X4 _35616_ (.A(_11665_),
    .ZN(_15313_));
 INV_X2 _35617_ (.A(_11655_),
    .ZN(_15155_));
 NOR2_X1 _35618_ (.A1(_15313_),
    .A2(_15155_),
    .ZN(_20649_));
 AND2_X1 _35619_ (.A1(_11642_),
    .A2(_11645_),
    .ZN(_14547_));
 AND2_X1 _35620_ (.A1(_11649_),
    .A2(_11654_),
    .ZN(_14546_));
 AND2_X1 _35621_ (.A1(_11644_),
    .A2(_11651_),
    .ZN(_14548_));
 AND2_X1 _35622_ (.A1(_11658_),
    .A2(_11663_),
    .ZN(_14551_));
 BUF_X1 _35623_ (.A(_11647_),
    .Z(_11666_));
 AND2_X1 _35624_ (.A1(_11666_),
    .A2(_11652_),
    .ZN(_14552_));
 AND2_X1 _35625_ (.A1(_11646_),
    .A2(_11660_),
    .ZN(_14553_));
 AND2_X1 _35626_ (.A1(_11646_),
    .A2(_11663_),
    .ZN(_20652_));
 AND2_X1 _35627_ (.A1(_11652_),
    .A2(_11660_),
    .ZN(_20653_));
 AND2_X1 _35628_ (.A1(_11666_),
    .A2(_11649_),
    .ZN(_14564_));
 AND2_X1 _35629_ (.A1(_11642_),
    .A2(_11651_),
    .ZN(_14565_));
 AND2_X1 _35630_ (.A1(_11644_),
    .A2(_11653_),
    .ZN(_14566_));
 BUF_X1 _35631_ (.A(net232),
    .Z(_11667_));
 BUF_X4 _35632_ (.A(_11667_),
    .Z(_11668_));
 AND2_X1 _35633_ (.A1(_11668_),
    .A2(_11655_),
    .ZN(_14596_));
 AND2_X1 _35634_ (.A1(_11664_),
    .A2(_11658_),
    .ZN(_14595_));
 BUF_X2 _35635_ (.A(_11665_),
    .Z(_11669_));
 AND2_X1 _35636_ (.A1(_11669_),
    .A2(_11661_),
    .ZN(_14594_));
 AND2_X1 _35637_ (.A1(_11642_),
    .A2(_11653_),
    .ZN(_20654_));
 AND2_X1 _35638_ (.A1(_11644_),
    .A2(_11648_),
    .ZN(_20655_));
 BUF_X1 _35639_ (.A(net267),
    .Z(_11670_));
 BUF_X1 _35640_ (.A(_11670_),
    .Z(_11671_));
 BUF_X2 _35641_ (.A(a[183]),
    .Z(_11672_));
 AND2_X1 _35642_ (.A1(_11671_),
    .A2(_11672_),
    .ZN(_14583_));
 BUF_X1 _35643_ (.A(b[57]),
    .Z(_11673_));
 CLKBUF_X3 _35644_ (.A(_11673_),
    .Z(_11674_));
 BUF_X2 _35645_ (.A(net83),
    .Z(_11675_));
 AND2_X1 _35646_ (.A1(_11674_),
    .A2(_11675_),
    .ZN(_14582_));
 INV_X1 _35647_ (.A(_11673_),
    .ZN(_18850_));
 INV_X2 _35648_ (.A(_11672_),
    .ZN(_14569_));
 NOR2_X1 _35649_ (.A1(_18850_),
    .A2(_14569_),
    .ZN(_14580_));
 BUF_X2 _35650_ (.A(net84),
    .Z(_11676_));
 BUF_X1 _35651_ (.A(net266),
    .Z(_11677_));
 BUF_X2 _35652_ (.A(_11677_),
    .Z(_11678_));
 AND2_X1 _35653_ (.A1(_11676_),
    .A2(_11678_),
    .ZN(_15322_));
 BUF_X2 _35654_ (.A(a[185]),
    .Z(_11679_));
 INV_X2 _35655_ (.A(_11679_),
    .ZN(_19209_));
 BUF_X2 _35656_ (.A(b[54]),
    .Z(_11680_));
 INV_X4 _35657_ (.A(_11680_),
    .ZN(_14944_));
 NOR2_X1 _35658_ (.A1(_19209_),
    .A2(_14944_),
    .ZN(_15323_));
 AND2_X1 _35659_ (.A1(_11671_),
    .A2(_11675_),
    .ZN(_15253_));
 BUF_X2 _35660_ (.A(net82),
    .Z(_11681_));
 AND2_X1 _35661_ (.A1(_11674_),
    .A2(_11681_),
    .ZN(_15252_));
 CLKBUF_X3 _35662_ (.A(_11677_),
    .Z(_11682_));
 AND2_X1 _35663_ (.A1(_11682_),
    .A2(_11672_),
    .ZN(_15247_));
 BUF_X1 _35664_ (.A(net265),
    .Z(_11683_));
 BUF_X1 _35665_ (.A(_11683_),
    .Z(_11684_));
 AND2_X1 _35666_ (.A1(_11679_),
    .A2(_11684_),
    .ZN(_15248_));
 AND2_X1 _35667_ (.A1(_11676_),
    .A2(_11680_),
    .ZN(_15249_));
 AND2_X1 _35668_ (.A1(_11646_),
    .A2(_11657_),
    .ZN(_14608_));
 AND2_X1 _35669_ (.A1(_11649_),
    .A2(_11660_),
    .ZN(_14609_));
 AND2_X1 _35670_ (.A1(_11652_),
    .A2(_11663_),
    .ZN(_14610_));
 AND2_X1 _35671_ (.A1(_11642_),
    .A2(_11648_),
    .ZN(_14625_));
 AND2_X1 _35672_ (.A1(_11649_),
    .A2(_11662_),
    .ZN(_14624_));
 AND2_X1 _35673_ (.A1(_11644_),
    .A2(_11660_),
    .ZN(_14626_));
 AND2_X1 _35674_ (.A1(_11652_),
    .A2(_11657_),
    .ZN(_20658_));
 AND2_X1 _35675_ (.A1(_11669_),
    .A2(_11646_),
    .ZN(_20659_));
 NOR2_X1 _35676_ (.A1(_19209_),
    .A2(_18850_),
    .ZN(_14613_));
 AND2_X1 _35677_ (.A1(_11644_),
    .A2(_11662_),
    .ZN(_20661_));
 AND2_X1 _35678_ (.A1(_11642_),
    .A2(_11660_),
    .ZN(_20662_));
 AND2_X1 _35679_ (.A1(_11668_),
    .A2(_11646_),
    .ZN(_14635_));
 AND2_X1 _35680_ (.A1(_11649_),
    .A2(_11657_),
    .ZN(_14634_));
 AND2_X1 _35681_ (.A1(_11669_),
    .A2(_11652_),
    .ZN(_14633_));
 BUF_X1 _35682_ (.A(net1),
    .Z(_11685_));
 AND2_X1 _35683_ (.A1(_11664_),
    .A2(_11685_),
    .ZN(_21086_));
 BUF_X2 _35684_ (.A(net100),
    .Z(_11686_));
 AND2_X1 _35685_ (.A1(_11669_),
    .A2(_11686_),
    .ZN(_21087_));
 AND2_X1 _35686_ (.A1(_11642_),
    .A2(_11662_),
    .ZN(_20664_));
 AND2_X1 _35687_ (.A1(_11644_),
    .A2(_11657_),
    .ZN(_20663_));
 AND2_X1 _35688_ (.A1(_11642_),
    .A2(_11657_),
    .ZN(_21102_));
 AND2_X1 _35689_ (.A1(_11669_),
    .A2(_11644_),
    .ZN(_21103_));
 BUF_X2 _35690_ (.A(net142),
    .Z(_11687_));
 BUF_X1 _35691_ (.A(b[49]),
    .Z(_11688_));
 AND2_X1 _35692_ (.A1(_11687_),
    .A2(_11688_),
    .ZN(_21117_));
 BUF_X2 _35693_ (.A(net141),
    .Z(_11689_));
 BUF_X1 _35694_ (.A(net263),
    .Z(_11690_));
 BUF_X1 _35695_ (.A(_11690_),
    .Z(_11691_));
 AND2_X1 _35696_ (.A1(_11689_),
    .A2(_11691_),
    .ZN(_21116_));
 CLKBUF_X3 _35697_ (.A(b[51]),
    .Z(_11692_));
 CLKBUF_X3 _35698_ (.A(_11692_),
    .Z(_11693_));
 AND2_X1 _35699_ (.A1(_11689_),
    .A2(_11693_),
    .ZN(_20667_));
 AND2_X1 _35700_ (.A1(_11687_),
    .A2(_11691_),
    .ZN(_20666_));
 BUF_X2 _35701_ (.A(a[167]),
    .Z(_11694_));
 INV_X2 _35702_ (.A(_11694_),
    .ZN(_16722_));
 CLKBUF_X3 _35703_ (.A(b[35]),
    .Z(_11695_));
 INV_X4 _35704_ (.A(_11695_),
    .ZN(_15412_));
 NOR2_X1 _35705_ (.A1(_16722_),
    .A2(_15412_),
    .ZN(_14647_));
 BUF_X2 _35706_ (.A(net66),
    .Z(_11696_));
 BUF_X1 _35707_ (.A(net253),
    .Z(_11697_));
 BUF_X1 _35708_ (.A(_11697_),
    .Z(_11698_));
 AND2_X1 _35709_ (.A1(_11696_),
    .A2(_11698_),
    .ZN(_14648_));
 BUF_X2 _35710_ (.A(net67),
    .Z(_11699_));
 BUF_X1 _35711_ (.A(net252),
    .Z(_11700_));
 CLKBUF_X3 _35712_ (.A(_11700_),
    .Z(_11701_));
 AND2_X1 _35713_ (.A1(_11699_),
    .A2(_11701_),
    .ZN(_14649_));
 BUF_X2 _35714_ (.A(net62),
    .Z(_11702_));
 BUF_X1 _35715_ (.A(net255),
    .Z(_11703_));
 AND2_X1 _35716_ (.A1(_11702_),
    .A2(_11703_),
    .ZN(_20673_));
 BUF_X2 _35717_ (.A(net64),
    .Z(_11704_));
 BUF_X1 _35718_ (.A(net254),
    .Z(_11705_));
 BUF_X2 _35719_ (.A(_11705_),
    .Z(_11706_));
 AND2_X1 _35720_ (.A1(_11704_),
    .A2(_11706_),
    .ZN(_20670_));
 BUF_X2 _35721_ (.A(net65),
    .Z(_11707_));
 CLKBUF_X3 _35722_ (.A(b[38]),
    .Z(_11708_));
 BUF_X2 _35723_ (.A(_11708_),
    .Z(_11709_));
 AND2_X1 _35724_ (.A1(_11707_),
    .A2(_11709_),
    .ZN(_20669_));
 BUF_X1 _35725_ (.A(_11703_),
    .Z(_11710_));
 BUF_X2 _35726_ (.A(net63),
    .Z(_11711_));
 AND2_X1 _35727_ (.A1(_11710_),
    .A2(_11711_),
    .ZN(_14638_));
 BUF_X1 _35728_ (.A(b[41]),
    .Z(_11712_));
 CLKBUF_X3 _35729_ (.A(_11712_),
    .Z(_11713_));
 AND2_X1 _35730_ (.A1(_11713_),
    .A2(_11702_),
    .ZN(_14639_));
 BUF_X2 _35731_ (.A(net68),
    .Z(_11714_));
 BUF_X1 _35732_ (.A(net251),
    .Z(_11715_));
 BUF_X1 _35733_ (.A(_11715_),
    .Z(_11716_));
 AND2_X1 _35734_ (.A1(_11714_),
    .A2(_11716_),
    .ZN(_14657_));
 BUF_X2 _35735_ (.A(a[169]),
    .Z(_11717_));
 INV_X2 _35736_ (.A(_11717_),
    .ZN(_19165_));
 BUF_X1 _35737_ (.A(b[33]),
    .Z(_11718_));
 INV_X4 _35738_ (.A(_11718_),
    .ZN(_14677_));
 NOR2_X1 _35739_ (.A1(_19165_),
    .A2(_14677_),
    .ZN(_14656_));
 BUF_X1 _35740_ (.A(_11697_),
    .Z(_11719_));
 AND2_X1 _35741_ (.A1(_11719_),
    .A2(_11707_),
    .ZN(_14690_));
 BUF_X4 _35742_ (.A(_11705_),
    .Z(_11720_));
 AND2_X1 _35743_ (.A1(_11720_),
    .A2(_11711_),
    .ZN(_14691_));
 AND2_X1 _35744_ (.A1(_11704_),
    .A2(_11709_),
    .ZN(_14692_));
 AND2_X1 _35745_ (.A1(_11696_),
    .A2(_11701_),
    .ZN(_14699_));
 AND2_X1 _35746_ (.A1(_11694_),
    .A2(_11716_),
    .ZN(_14700_));
 BUF_X2 _35747_ (.A(_11695_),
    .Z(_11721_));
 AND2_X1 _35748_ (.A1(_11721_),
    .A2(_11699_),
    .ZN(_14701_));
 AND2_X1 _35749_ (.A1(_11721_),
    .A2(_11714_),
    .ZN(_14666_));
 AND2_X1 _35750_ (.A1(_11719_),
    .A2(_11699_),
    .ZN(_14665_));
 AND2_X1 _35751_ (.A1(_11694_),
    .A2(_11701_),
    .ZN(_14664_));
 AND2_X1 _35752_ (.A1(_11696_),
    .A2(_11708_),
    .ZN(_20677_));
 AND2_X1 _35753_ (.A1(_11720_),
    .A2(_11707_),
    .ZN(_20676_));
 AND2_X1 _35754_ (.A1(_11710_),
    .A2(_11704_),
    .ZN(_14669_));
 AND2_X1 _35755_ (.A1(_11713_),
    .A2(_11711_),
    .ZN(_14670_));
 AND2_X1 _35756_ (.A1(_11699_),
    .A2(_11716_),
    .ZN(_20888_));
 NOR2_X1 _35757_ (.A1(_16722_),
    .A2(_14677_),
    .ZN(_20889_));
 BUF_X1 _35758_ (.A(net61),
    .Z(_11722_));
 AND2_X1 _35759_ (.A1(_11722_),
    .A2(_11703_),
    .ZN(_16704_));
 BUF_X2 _35760_ (.A(_11708_),
    .Z(_11723_));
 AND2_X1 _35761_ (.A1(_11723_),
    .A2(_11711_),
    .ZN(_16703_));
 AND2_X1 _35762_ (.A1(_11702_),
    .A2(_11706_),
    .ZN(_16702_));
 AND2_X1 _35763_ (.A1(_11719_),
    .A2(_11704_),
    .ZN(_16706_));
 AND2_X1 _35764_ (.A1(_11721_),
    .A2(_11696_),
    .ZN(_16707_));
 BUF_X1 _35765_ (.A(_11700_),
    .Z(_11724_));
 AND2_X1 _35766_ (.A1(_11724_),
    .A2(_11707_),
    .ZN(_16708_));
 AND2_X1 _35767_ (.A1(_11687_),
    .A2(_11693_),
    .ZN(_20679_));
 BUF_X1 _35768_ (.A(net264),
    .Z(_11725_));
 CLKBUF_X3 _35769_ (.A(_11725_),
    .Z(_11726_));
 AND2_X1 _35770_ (.A1(_11689_),
    .A2(_11726_),
    .ZN(_20678_));
 BUF_X1 _35771_ (.A(net261),
    .Z(_11727_));
 BUF_X4 _35772_ (.A(_11727_),
    .Z(_11728_));
 BUF_X2 _35773_ (.A(net145),
    .Z(_11729_));
 AND2_X1 _35774_ (.A1(_11728_),
    .A2(_11729_),
    .ZN(_14705_));
 BUF_X1 _35775_ (.A(_11690_),
    .Z(_11730_));
 BUF_X2 _35776_ (.A(net143),
    .Z(_11731_));
 AND2_X1 _35777_ (.A1(_11730_),
    .A2(_11731_),
    .ZN(_14704_));
 BUF_X1 _35778_ (.A(_11688_),
    .Z(_11732_));
 BUF_X2 _35779_ (.A(net144),
    .Z(_11733_));
 AND2_X1 _35780_ (.A1(_11732_),
    .A2(_11733_),
    .ZN(_14706_));
 AND2_X1 _35781_ (.A1(_11730_),
    .A2(_11733_),
    .ZN(_20681_));
 AND2_X1 _35782_ (.A1(_11732_),
    .A2(_11729_),
    .ZN(_20682_));
 BUF_X1 _35783_ (.A(_11683_),
    .Z(_11734_));
 AND2_X1 _35784_ (.A1(_11734_),
    .A2(_11689_),
    .ZN(_14711_));
 AND2_X1 _35785_ (.A1(_11731_),
    .A2(_11693_),
    .ZN(_14710_));
 AND2_X1 _35786_ (.A1(_11687_),
    .A2(_11726_),
    .ZN(_14709_));
 BUF_X2 _35787_ (.A(_11680_),
    .Z(_11735_));
 AND2_X1 _35788_ (.A1(_11735_),
    .A2(_11689_),
    .ZN(_20684_));
 AND2_X1 _35789_ (.A1(_11734_),
    .A2(_11687_),
    .ZN(_20683_));
 AND2_X1 _35790_ (.A1(_11730_),
    .A2(_11729_),
    .ZN(_14724_));
 AND2_X1 _35791_ (.A1(_11731_),
    .A2(_11726_),
    .ZN(_14725_));
 BUF_X2 _35792_ (.A(_11692_),
    .Z(_11736_));
 AND2_X1 _35793_ (.A1(_11736_),
    .A2(_11733_),
    .ZN(_14726_));
 AND2_X1 _35794_ (.A1(_11736_),
    .A2(_11729_),
    .ZN(_20686_));
 AND2_X1 _35795_ (.A1(_11733_),
    .A2(_11726_),
    .ZN(_20687_));
 AND2_X1 _35796_ (.A1(_11734_),
    .A2(_11731_),
    .ZN(_14732_));
 AND2_X1 _35797_ (.A1(_11682_),
    .A2(_11689_),
    .ZN(_14733_));
 AND2_X1 _35798_ (.A1(_11735_),
    .A2(_11687_),
    .ZN(_14734_));
 BUF_X2 _35799_ (.A(a[247]),
    .Z(_11737_));
 AND2_X1 _35800_ (.A1(_11728_),
    .A2(_11737_),
    .ZN(_14742_));
 BUF_X2 _35801_ (.A(net146),
    .Z(_11738_));
 AND2_X1 _35802_ (.A1(_11730_),
    .A2(_11738_),
    .ZN(_14741_));
 BUF_X2 _35803_ (.A(net147),
    .Z(_11739_));
 AND2_X1 _35804_ (.A1(_11732_),
    .A2(_11739_),
    .ZN(_14743_));
 AND2_X1 _35805_ (.A1(_11671_),
    .A2(_11689_),
    .ZN(_14750_));
 AND2_X1 _35806_ (.A1(_11735_),
    .A2(_11731_),
    .ZN(_14751_));
 AND2_X1 _35807_ (.A1(_11682_),
    .A2(_11687_),
    .ZN(_14752_));
 AND2_X1 _35808_ (.A1(_11730_),
    .A2(_11739_),
    .ZN(_20690_));
 INV_X4 _35809_ (.A(_11688_),
    .ZN(_14841_));
 INV_X2 _35810_ (.A(_11737_),
    .ZN(_14957_));
 NOR2_X1 _35811_ (.A1(_14841_),
    .A2(_14957_),
    .ZN(_20689_));
 AND2_X1 _35812_ (.A1(_11736_),
    .A2(_11738_),
    .ZN(_14757_));
 AND2_X1 _35813_ (.A1(_11734_),
    .A2(_11733_),
    .ZN(_14756_));
 CLKBUF_X3 _35814_ (.A(_11725_),
    .Z(_11740_));
 AND2_X1 _35815_ (.A1(_11740_),
    .A2(_11729_),
    .ZN(_14755_));
 AND2_X1 _35816_ (.A1(_11682_),
    .A2(_11731_),
    .ZN(_14776_));
 AND2_X1 _35817_ (.A1(_11734_),
    .A2(_11729_),
    .ZN(_14775_));
 AND2_X1 _35818_ (.A1(_11735_),
    .A2(_11733_),
    .ZN(_14774_));
 AND2_X1 _35819_ (.A1(_11674_),
    .A2(_11689_),
    .ZN(_20692_));
 AND2_X1 _35820_ (.A1(_11671_),
    .A2(_11687_),
    .ZN(_20693_));
 AND2_X1 _35821_ (.A1(_11730_),
    .A2(_11737_),
    .ZN(_14786_));
 AND2_X1 _35822_ (.A1(_11740_),
    .A2(_11738_),
    .ZN(_14785_));
 AND2_X1 _35823_ (.A1(_11736_),
    .A2(_11739_),
    .ZN(_14784_));
 AND2_X1 _35824_ (.A1(_11682_),
    .A2(_11733_),
    .ZN(_20695_));
 AND2_X1 _35825_ (.A1(_11735_),
    .A2(_11729_),
    .ZN(_20696_));
 AND2_X1 _35826_ (.A1(_11671_),
    .A2(_11731_),
    .ZN(_14800_));
 AND2_X1 _35827_ (.A1(_11674_),
    .A2(_11687_),
    .ZN(_14799_));
 AND2_X1 _35828_ (.A1(_11734_),
    .A2(_11738_),
    .ZN(_14807_));
 INV_X4 _35829_ (.A(_11692_),
    .ZN(_14888_));
 NOR2_X1 _35830_ (.A1(_14888_),
    .A2(_14957_),
    .ZN(_14808_));
 AND2_X1 _35831_ (.A1(_11740_),
    .A2(_11739_),
    .ZN(_14809_));
 BUF_X1 _35832_ (.A(_11690_),
    .Z(_11741_));
 BUF_X2 _35833_ (.A(net148),
    .Z(_11742_));
 AND2_X1 _35834_ (.A1(_11741_),
    .A2(_11742_),
    .ZN(_14813_));
 BUF_X2 _35835_ (.A(a[249]),
    .Z(_11743_));
 INV_X2 _35836_ (.A(_11743_),
    .ZN(_19397_));
 NOR2_X1 _35837_ (.A1(_14841_),
    .A2(_19397_),
    .ZN(_14812_));
 AND2_X1 _35838_ (.A1(_11682_),
    .A2(_11729_),
    .ZN(_20698_));
 AND2_X1 _35839_ (.A1(_11735_),
    .A2(_11738_),
    .ZN(_20697_));
 AND2_X1 _35840_ (.A1(_11671_),
    .A2(_11733_),
    .ZN(_14828_));
 AND2_X1 _35841_ (.A1(_11674_),
    .A2(_11731_),
    .ZN(_14829_));
 AND2_X1 _35842_ (.A1(_11736_),
    .A2(_11742_),
    .ZN(_14838_));
 AND2_X1 _35843_ (.A1(_11734_),
    .A2(_11739_),
    .ZN(_14837_));
 AND2_X1 _35844_ (.A1(_11740_),
    .A2(_11737_),
    .ZN(_14836_));
 BUF_X2 _35845_ (.A(_11677_),
    .Z(_11744_));
 AND2_X1 _35846_ (.A1(_11744_),
    .A2(_11738_),
    .ZN(_14857_));
 AND2_X1 _35847_ (.A1(_11734_),
    .A2(_11737_),
    .ZN(_14858_));
 AND2_X1 _35848_ (.A1(_11735_),
    .A2(_11739_),
    .ZN(_14859_));
 BUF_X1 _35849_ (.A(_11670_),
    .Z(_11745_));
 AND2_X1 _35850_ (.A1(_11745_),
    .A2(_11729_),
    .ZN(_14863_));
 AND2_X1 _35851_ (.A1(_11674_),
    .A2(_11733_),
    .ZN(_14862_));
 AND2_X1 _35852_ (.A1(_11740_),
    .A2(_11742_),
    .ZN(_14869_));
 NOR2_X1 _35853_ (.A1(_14888_),
    .A2(_19397_),
    .ZN(_14870_));
 AND2_X1 _35854_ (.A1(_11745_),
    .A2(_11738_),
    .ZN(_14884_));
 BUF_X2 _35855_ (.A(_11673_),
    .Z(_11746_));
 AND2_X1 _35856_ (.A1(_11746_),
    .A2(_11729_),
    .ZN(_14885_));
 AND2_X1 _35857_ (.A1(_11744_),
    .A2(_11739_),
    .ZN(_14893_));
 AND2_X1 _35858_ (.A1(_11734_),
    .A2(_11742_),
    .ZN(_14894_));
 NOR2_X1 _35859_ (.A1(_14944_),
    .A2(_14957_),
    .ZN(_14895_));
 AND2_X1 _35860_ (.A1(_11734_),
    .A2(_11743_),
    .ZN(_14909_));
 AND2_X1 _35861_ (.A1(_11744_),
    .A2(_11737_),
    .ZN(_14910_));
 AND2_X1 _35862_ (.A1(_11735_),
    .A2(_11742_),
    .ZN(_14911_));
 AND2_X1 _35863_ (.A1(_11745_),
    .A2(_11739_),
    .ZN(_14914_));
 AND2_X1 _35864_ (.A1(_11746_),
    .A2(_11738_),
    .ZN(_14915_));
 AND2_X1 _35865_ (.A1(_11745_),
    .A2(_11737_),
    .ZN(_14927_));
 AND2_X1 _35866_ (.A1(_11746_),
    .A2(_11739_),
    .ZN(_14928_));
 AND2_X1 _35867_ (.A1(_11744_),
    .A2(_11742_),
    .ZN(_14937_));
 NOR2_X1 _35868_ (.A1(_14944_),
    .A2(_19397_),
    .ZN(_14936_));
 NOR2_X1 _35869_ (.A1(_18850_),
    .A2(_14957_),
    .ZN(_14950_));
 NOR2_X1 _35870_ (.A1(_18850_),
    .A2(_19397_),
    .ZN(_14965_));
 INV_X4 _35871_ (.A(_11662_),
    .ZN(_15238_));
 NOR2_X1 _35872_ (.A1(_15155_),
    .A2(_15238_),
    .ZN(_14968_));
 AND2_X1 _35873_ (.A1(_11666_),
    .A2(_11658_),
    .ZN(_14969_));
 CLKBUF_X3 _35874_ (.A(_11659_),
    .Z(_11747_));
 AND2_X1 _35875_ (.A1(_11747_),
    .A2(_11661_),
    .ZN(_14970_));
 CLKBUF_X3 _35876_ (.A(_11650_),
    .Z(_11748_));
 AND2_X1 _35877_ (.A1(_11748_),
    .A2(_11652_),
    .ZN(_20701_));
 AND2_X1 _35878_ (.A1(_11646_),
    .A2(_11653_),
    .ZN(_20700_));
 BUF_X1 _35879_ (.A(_11645_),
    .Z(_11749_));
 AND2_X1 _35880_ (.A1(_11749_),
    .A2(_11649_),
    .ZN(_14973_));
 CLKBUF_X3 _35881_ (.A(_11643_),
    .Z(_11750_));
 AND2_X1 _35882_ (.A1(_11750_),
    .A2(_11644_),
    .ZN(_14974_));
 BUF_X2 _35883_ (.A(net36),
    .Z(_11751_));
 AND2_X1 _35884_ (.A1(_11751_),
    .A2(_11657_),
    .ZN(_14982_));
 BUF_X2 _35885_ (.A(a[137]),
    .Z(_11752_));
 INV_X2 _35886_ (.A(_11752_),
    .ZN(_19072_));
 NOR2_X1 _35887_ (.A1(_15313_),
    .A2(_19072_),
    .ZN(_14981_));
 BUF_X2 _35888_ (.A(net78),
    .Z(_11753_));
 AND2_X1 _35889_ (.A1(_11735_),
    .A2(_11753_),
    .ZN(_15002_));
 BUF_X2 _35890_ (.A(net76),
    .Z(_11754_));
 AND2_X1 _35891_ (.A1(_11745_),
    .A2(_11754_),
    .ZN(_15003_));
 BUF_X2 _35892_ (.A(net77),
    .Z(_11755_));
 AND2_X1 _35893_ (.A1(_11744_),
    .A2(_11755_),
    .ZN(_15001_));
 AND2_X1 _35894_ (.A1(_11675_),
    .A2(_11691_),
    .ZN(_20705_));
 NOR2_X1 _35895_ (.A1(_14569_),
    .A2(_14841_),
    .ZN(_20704_));
 BUF_X1 _35896_ (.A(_11683_),
    .Z(_11756_));
 BUF_X2 _35897_ (.A(net79),
    .Z(_11757_));
 AND2_X1 _35898_ (.A1(_11756_),
    .A2(_11757_),
    .ZN(_15005_));
 AND2_X1 _35899_ (.A1(_11681_),
    .A2(_11693_),
    .ZN(_15006_));
 BUF_X2 _35900_ (.A(net81),
    .Z(_11758_));
 AND2_X1 _35901_ (.A1(_11740_),
    .A2(_11758_),
    .ZN(_15007_));
 BUF_X2 _35902_ (.A(_11725_),
    .Z(_11759_));
 AND2_X1 _35903_ (.A1(_11759_),
    .A2(_11757_),
    .ZN(_20712_));
 AND2_X1 _35904_ (.A1(_11736_),
    .A2(_11758_),
    .ZN(_20711_));
 AND2_X1 _35905_ (.A1(_11756_),
    .A2(_11753_),
    .ZN(_15037_));
 AND2_X1 _35906_ (.A1(_11744_),
    .A2(_11754_),
    .ZN(_15038_));
 AND2_X1 _35907_ (.A1(_11735_),
    .A2(_11755_),
    .ZN(_15039_));
 AND2_X1 _35908_ (.A1(_11756_),
    .A2(_11758_),
    .ZN(_15014_));
 AND2_X1 _35909_ (.A1(_11744_),
    .A2(_11753_),
    .ZN(_15015_));
 BUF_X2 _35910_ (.A(_11680_),
    .Z(_11760_));
 AND2_X1 _35911_ (.A1(_11760_),
    .A2(_11757_),
    .ZN(_15016_));
 AND2_X1 _35912_ (.A1(_11745_),
    .A2(_11755_),
    .ZN(_20707_));
 AND2_X1 _35913_ (.A1(_11681_),
    .A2(_11726_),
    .ZN(_15024_));
 AND2_X1 _35914_ (.A1(_11672_),
    .A2(_11691_),
    .ZN(_15025_));
 AND2_X1 _35915_ (.A1(_11675_),
    .A2(_11692_),
    .ZN(_15026_));
 AND2_X1 _35916_ (.A1(_11681_),
    .A2(_11691_),
    .ZN(_15665_));
 BUF_X1 _35917_ (.A(_11727_),
    .Z(_11761_));
 AND2_X1 _35918_ (.A1(_11672_),
    .A2(_11761_),
    .ZN(_15664_));
 AND2_X1 _35919_ (.A1(_11675_),
    .A2(_11688_),
    .ZN(_15663_));
 AND2_X1 _35920_ (.A1(_11760_),
    .A2(_11754_),
    .ZN(_20763_));
 BUF_X1 _35921_ (.A(net239),
    .Z(_11762_));
 BUF_X1 _35922_ (.A(_11762_),
    .Z(_11763_));
 BUF_X1 _35923_ (.A(net69),
    .Z(_11764_));
 AND2_X1 _35924_ (.A1(_11763_),
    .A2(_11764_),
    .ZN(_21088_));
 BUF_X4 _35925_ (.A(b[17]),
    .Z(_11765_));
 BUF_X4 _35926_ (.A(_11765_),
    .Z(_11766_));
 BUF_X2 _35927_ (.A(net80),
    .Z(_11767_));
 AND2_X1 _35928_ (.A1(_11766_),
    .A2(_11767_),
    .ZN(_21089_));
 NOR2_X1 _35929_ (.A1(_14569_),
    .A2(_14888_),
    .ZN(_15051_));
 AND2_X1 _35930_ (.A1(_11681_),
    .A2(_11684_),
    .ZN(_15050_));
 AND2_X1 _35931_ (.A1(_11675_),
    .A2(_11726_),
    .ZN(_15049_));
 AND2_X1 _35932_ (.A1(_11760_),
    .A2(_11758_),
    .ZN(_20715_));
 AND2_X1 _35933_ (.A1(_11744_),
    .A2(_11757_),
    .ZN(_20716_));
 AND2_X1 _35934_ (.A1(_11745_),
    .A2(_11753_),
    .ZN(_15054_));
 AND2_X1 _35935_ (.A1(_11746_),
    .A2(_11755_),
    .ZN(_15055_));
 AND2_X1 _35936_ (.A1(_11676_),
    .A2(_11691_),
    .ZN(_15064_));
 NOR2_X1 _35937_ (.A1(_19209_),
    .A2(_14841_),
    .ZN(_15063_));
 AND2_X1 _35938_ (.A1(_11760_),
    .A2(_11681_),
    .ZN(_20719_));
 AND2_X1 _35939_ (.A1(_11744_),
    .A2(_11758_),
    .ZN(_20718_));
 AND2_X1 _35940_ (.A1(_11745_),
    .A2(_11757_),
    .ZN(_15077_));
 AND2_X1 _35941_ (.A1(_11746_),
    .A2(_11753_),
    .ZN(_15078_));
 AND2_X1 _35942_ (.A1(_11675_),
    .A2(_11684_),
    .ZN(_15085_));
 AND2_X1 _35943_ (.A1(_11676_),
    .A2(_11692_),
    .ZN(_15086_));
 AND2_X1 _35944_ (.A1(_11672_),
    .A2(_11726_),
    .ZN(_15087_));
 INV_X1 _35945_ (.A(_11643_),
    .ZN(_18713_));
 NOR2_X1 _35946_ (.A1(_18713_),
    .A2(_19072_),
    .ZN(_15125_));
 AND2_X1 _35947_ (.A1(_11745_),
    .A2(_11758_),
    .ZN(_15104_));
 AND2_X1 _35948_ (.A1(_11746_),
    .A2(_11757_),
    .ZN(_15105_));
 AND2_X1 _35949_ (.A1(_11672_),
    .A2(_11684_),
    .ZN(_15111_));
 AND2_X1 _35950_ (.A1(_11744_),
    .A2(_11681_),
    .ZN(_15112_));
 AND2_X1 _35951_ (.A1(_11675_),
    .A2(_11680_),
    .ZN(_15113_));
 AND2_X1 _35952_ (.A1(_11676_),
    .A2(_11726_),
    .ZN(_15116_));
 NOR2_X1 _35953_ (.A1(_19209_),
    .A2(_14888_),
    .ZN(_15117_));
 AND2_X1 _35954_ (.A1(_11749_),
    .A2(_11655_),
    .ZN(_15169_));
 AND2_X1 _35955_ (.A1(_11750_),
    .A2(_11661_),
    .ZN(_15168_));
 NOR2_X1 _35956_ (.A1(_18713_),
    .A2(_15155_),
    .ZN(_15166_));
 AND2_X1 _35957_ (.A1(_11696_),
    .A2(_11706_),
    .ZN(_15134_));
 AND2_X1 _35958_ (.A1(_11694_),
    .A2(_11698_),
    .ZN(_15136_));
 AND2_X1 _35959_ (.A1(_11699_),
    .A2(_11708_),
    .ZN(_15135_));
 AND2_X1 _35960_ (.A1(_11710_),
    .A2(_11707_),
    .ZN(_15140_));
 AND2_X1 _35961_ (.A1(_11713_),
    .A2(_11704_),
    .ZN(_15139_));
 AND2_X1 _35962_ (.A1(_11724_),
    .A2(_11714_),
    .ZN(_15147_));
 NOR2_X1 _35963_ (.A1(_15412_),
    .A2(_19165_),
    .ZN(_15146_));
 AND2_X1 _35964_ (.A1(_11751_),
    .A2(_11651_),
    .ZN(_15206_));
 INV_X4 _35965_ (.A(_11653_),
    .ZN(_15196_));
 NOR2_X1 _35966_ (.A1(_19072_),
    .A2(_15196_),
    .ZN(_15205_));
 AND2_X1 _35967_ (.A1(_11749_),
    .A2(_11661_),
    .ZN(_15214_));
 AND2_X1 _35968_ (.A1(_11750_),
    .A2(_11658_),
    .ZN(_15215_));
 AND2_X1 _35969_ (.A1(_11748_),
    .A2(_11655_),
    .ZN(_15210_));
 AND2_X1 _35970_ (.A1(_11752_),
    .A2(_11648_),
    .ZN(_15209_));
 AND2_X1 _35971_ (.A1(_11751_),
    .A2(_11653_),
    .ZN(_15211_));
 AND2_X1 _35972_ (.A1(_11745_),
    .A2(_11681_),
    .ZN(_15173_));
 AND2_X1 _35973_ (.A1(_11746_),
    .A2(_11758_),
    .ZN(_15172_));
 AND2_X1 _35974_ (.A1(_11676_),
    .A2(_11684_),
    .ZN(_15180_));
 BUF_X2 _35975_ (.A(_11677_),
    .Z(_11768_));
 AND2_X1 _35976_ (.A1(_11768_),
    .A2(_11675_),
    .ZN(_15181_));
 NOR2_X1 _35977_ (.A1(_14569_),
    .A2(_14944_),
    .ZN(_15182_));
 AND2_X1 _35978_ (.A1(_11748_),
    .A2(_11661_),
    .ZN(_15244_));
 AND2_X1 _35979_ (.A1(_11751_),
    .A2(_11648_),
    .ZN(_15243_));
 NOR2_X1 _35980_ (.A1(_15196_),
    .A2(_15155_),
    .ZN(_15245_));
 AND2_X1 _35981_ (.A1(_11749_),
    .A2(_11658_),
    .ZN(_15235_));
 AND2_X1 _35982_ (.A1(_11750_),
    .A2(_11646_),
    .ZN(_15236_));
 AND2_X1 _35983_ (.A1(_11749_),
    .A2(_11646_),
    .ZN(_15227_));
 AND2_X1 _35984_ (.A1(_11750_),
    .A2(_11652_),
    .ZN(_15228_));
 AND2_X1 _35985_ (.A1(_11749_),
    .A2(_11652_),
    .ZN(_15277_));
 AND2_X1 _35986_ (.A1(_11750_),
    .A2(_11649_),
    .ZN(_15278_));
 AND2_X1 _35987_ (.A1(_11646_),
    .A2(_11651_),
    .ZN(_20721_));
 BUF_X2 _35988_ (.A(_11653_),
    .Z(_11769_));
 AND2_X1 _35989_ (.A1(_11769_),
    .A2(_11658_),
    .ZN(_20722_));
 AND2_X1 _35990_ (.A1(_11748_),
    .A2(_11658_),
    .ZN(_15282_));
 AND2_X1 _35991_ (.A1(_11666_),
    .A2(_11655_),
    .ZN(_15281_));
 AND2_X1 _35992_ (.A1(_11769_),
    .A2(_11661_),
    .ZN(_15283_));
 AND2_X1 _35993_ (.A1(_11751_),
    .A2(_11660_),
    .ZN(_15290_));
 NOR2_X1 _35994_ (.A1(_19072_),
    .A2(_15238_),
    .ZN(_15289_));
 AND2_X1 _35995_ (.A1(_11666_),
    .A2(_11661_),
    .ZN(_15304_));
 AND2_X1 _35996_ (.A1(_11751_),
    .A2(_11662_),
    .ZN(_15305_));
 AND2_X1 _35997_ (.A1(_11655_),
    .A2(_11660_),
    .ZN(_15306_));
 AND2_X1 _35998_ (.A1(_11741_),
    .A2(_11754_),
    .ZN(_21109_));
 AND2_X1 _35999_ (.A1(_11732_),
    .A2(_11755_),
    .ZN(_21108_));
 BUF_X1 _36000_ (.A(_11715_),
    .Z(_11770_));
 BUF_X2 _36001_ (.A(net163),
    .Z(_11771_));
 AND2_X1 _36002_ (.A1(_11770_),
    .A2(_11771_),
    .ZN(_21091_));
 BUF_X1 _36003_ (.A(_11718_),
    .Z(_11772_));
 BUF_X2 _36004_ (.A(net164),
    .Z(_11773_));
 AND2_X1 _36005_ (.A1(_11772_),
    .A2(_11773_),
    .ZN(_21090_));
 AND2_X1 _36006_ (.A1(_11741_),
    .A2(_11755_),
    .ZN(_20725_));
 AND2_X1 _36007_ (.A1(_11736_),
    .A2(_11754_),
    .ZN(_20724_));
 BUF_X2 _36008_ (.A(net125),
    .Z(_11774_));
 AND2_X1 _36009_ (.A1(_11770_),
    .A2(_11774_),
    .ZN(_21114_));
 BUF_X2 _36010_ (.A(net126),
    .Z(_11775_));
 AND2_X1 _36011_ (.A1(_11772_),
    .A2(_11775_),
    .ZN(_21115_));
 AND2_X1 _36012_ (.A1(_11721_),
    .A2(_11774_),
    .ZN(_20727_));
 AND2_X1 _36013_ (.A1(_11770_),
    .A2(_11775_),
    .ZN(_20728_));
 BUF_X1 _36014_ (.A(net250),
    .Z(_11776_));
 BUF_X4 _36015_ (.A(_11776_),
    .Z(_11777_));
 BUF_X2 _36016_ (.A(net129),
    .Z(_11778_));
 AND2_X1 _36017_ (.A1(_11777_),
    .A2(_11778_),
    .ZN(_15355_));
 BUF_X2 _36018_ (.A(net127),
    .Z(_11779_));
 AND2_X1 _36019_ (.A1(_11770_),
    .A2(_11779_),
    .ZN(_15354_));
 BUF_X2 _36020_ (.A(net128),
    .Z(_11780_));
 AND2_X1 _36021_ (.A1(_11772_),
    .A2(_11780_),
    .ZN(_15353_));
 AND2_X1 _36022_ (.A1(_11724_),
    .A2(_11774_),
    .ZN(_20730_));
 AND2_X1 _36023_ (.A1(_11721_),
    .A2(_11775_),
    .ZN(_20731_));
 AND2_X1 _36024_ (.A1(_11721_),
    .A2(_11779_),
    .ZN(_15358_));
 AND2_X1 _36025_ (.A1(_11719_),
    .A2(_11774_),
    .ZN(_15359_));
 AND2_X1 _36026_ (.A1(_11724_),
    .A2(_11775_),
    .ZN(_15360_));
 AND2_X1 _36027_ (.A1(_11770_),
    .A2(_11780_),
    .ZN(_20733_));
 AND2_X1 _36028_ (.A1(_11772_),
    .A2(_11778_),
    .ZN(_20734_));
 BUF_X1 _36029_ (.A(_11727_),
    .Z(_11781_));
 AND2_X1 _36030_ (.A1(_11781_),
    .A2(_11758_),
    .ZN(_15370_));
 AND2_X1 _36031_ (.A1(_11741_),
    .A2(_11753_),
    .ZN(_15369_));
 AND2_X1 _36032_ (.A1(_11732_),
    .A2(_11757_),
    .ZN(_15368_));
 AND2_X1 _36033_ (.A1(_11759_),
    .A2(_11754_),
    .ZN(_20736_));
 AND2_X1 _36034_ (.A1(_11736_),
    .A2(_11755_),
    .ZN(_20737_));
 AND2_X1 _36035_ (.A1(_11770_),
    .A2(_11778_),
    .ZN(_15373_));
 AND2_X1 _36036_ (.A1(_11724_),
    .A2(_11779_),
    .ZN(_15374_));
 AND2_X1 _36037_ (.A1(_11721_),
    .A2(_11780_),
    .ZN(_15375_));
 AND2_X1 _36038_ (.A1(_11723_),
    .A2(_11774_),
    .ZN(_20739_));
 BUF_X2 _36039_ (.A(_11715_),
    .Z(_11782_));
 BUF_X2 _36040_ (.A(net130),
    .Z(_11783_));
 AND2_X1 _36041_ (.A1(_11782_),
    .A2(_11783_),
    .ZN(_15386_));
 BUF_X2 _36042_ (.A(net133),
    .Z(_11784_));
 AND2_X1 _36043_ (.A1(_11777_),
    .A2(_11784_),
    .ZN(_15388_));
 BUF_X2 _36044_ (.A(net132),
    .Z(_11785_));
 AND2_X1 _36045_ (.A1(_11772_),
    .A2(_11785_),
    .ZN(_15387_));
 AND2_X1 _36046_ (.A1(_11724_),
    .A2(_11780_),
    .ZN(_20743_));
 AND2_X1 _36047_ (.A1(_11721_),
    .A2(_11778_),
    .ZN(_20744_));
 AND2_X1 _36048_ (.A1(_11720_),
    .A2(_11774_),
    .ZN(_15395_));
 AND2_X1 _36049_ (.A1(_11719_),
    .A2(_11779_),
    .ZN(_15396_));
 AND2_X1 _36050_ (.A1(_11723_),
    .A2(_11775_),
    .ZN(_15397_));
 AND2_X1 _36051_ (.A1(_11696_),
    .A2(_11703_),
    .ZN(_15418_));
 AND2_X1 _36052_ (.A1(_11713_),
    .A2(_11707_),
    .ZN(_15417_));
 AND2_X1 _36053_ (.A1(_11719_),
    .A2(_11714_),
    .ZN(_15421_));
 AND2_X1 _36054_ (.A1(_11699_),
    .A2(_11706_),
    .ZN(_15422_));
 INV_X4 _36055_ (.A(_11708_),
    .ZN(_15651_));
 NOR2_X1 _36056_ (.A1(_16722_),
    .A2(_15651_),
    .ZN(_15423_));
 AND2_X1 _36057_ (.A1(_11782_),
    .A2(_11785_),
    .ZN(_20747_));
 AND2_X1 _36058_ (.A1(_11772_),
    .A2(_11784_),
    .ZN(_20748_));
 AND2_X1 _36059_ (.A1(_11723_),
    .A2(_11779_),
    .ZN(_15438_));
 AND2_X1 _36060_ (.A1(_11710_),
    .A2(_11774_),
    .ZN(_15439_));
 AND2_X1 _36061_ (.A1(_11720_),
    .A2(_11775_),
    .ZN(_15440_));
 AND2_X1 _36062_ (.A1(_11721_),
    .A2(_11783_),
    .ZN(_15443_));
 AND2_X1 _36063_ (.A1(_11719_),
    .A2(_11780_),
    .ZN(_15444_));
 CLKBUF_X3 _36064_ (.A(_11700_),
    .Z(_11786_));
 AND2_X1 _36065_ (.A1(_11786_),
    .A2(_11778_),
    .ZN(_15445_));
 AND2_X1 _36066_ (.A1(_11710_),
    .A2(_11775_),
    .ZN(_20750_));
 AND2_X1 _36067_ (.A1(_11720_),
    .A2(_11779_),
    .ZN(_15464_));
 AND2_X1 _36068_ (.A1(_11719_),
    .A2(_11778_),
    .ZN(_15465_));
 AND2_X1 _36069_ (.A1(_11723_),
    .A2(_11780_),
    .ZN(_15466_));
 AND2_X1 _36070_ (.A1(_11782_),
    .A2(_11784_),
    .ZN(_15471_));
 AND2_X1 _36071_ (.A1(_11786_),
    .A2(_11783_),
    .ZN(_15470_));
 AND2_X1 _36072_ (.A1(_11721_),
    .A2(_11785_),
    .ZN(_15469_));
 AND2_X1 _36073_ (.A1(_11756_),
    .A2(_11754_),
    .ZN(_15478_));
 AND2_X1 _36074_ (.A1(_11736_),
    .A2(_11753_),
    .ZN(_15479_));
 AND2_X1 _36075_ (.A1(_11759_),
    .A2(_11755_),
    .ZN(_15480_));
 AND2_X1 _36076_ (.A1(_11732_),
    .A2(_11758_),
    .ZN(_20755_));
 AND2_X1 _36077_ (.A1(_11741_),
    .A2(_11757_),
    .ZN(_20754_));
 CLKBUF_X3 _36078_ (.A(_11695_),
    .Z(_11787_));
 AND2_X1 _36079_ (.A1(_11787_),
    .A2(_11784_),
    .ZN(_15497_));
 AND2_X1 _36080_ (.A1(_11719_),
    .A2(_11783_),
    .ZN(_15496_));
 AND2_X1 _36081_ (.A1(_11786_),
    .A2(_11785_),
    .ZN(_15495_));
 AND2_X1 _36082_ (.A1(_11720_),
    .A2(_11780_),
    .ZN(_20757_));
 AND2_X1 _36083_ (.A1(_11723_),
    .A2(_11778_),
    .ZN(_20758_));
 AND2_X1 _36084_ (.A1(_11710_),
    .A2(_11779_),
    .ZN(_15500_));
 AND2_X1 _36085_ (.A1(_11713_),
    .A2(_11775_),
    .ZN(_15501_));
 BUF_X2 _36086_ (.A(net134),
    .Z(_11788_));
 AND2_X1 _36087_ (.A1(_11782_),
    .A2(_11788_),
    .ZN(_15510_));
 BUF_X2 _36088_ (.A(net352),
    .Z(_11789_));
 INV_X2 _36089_ (.A(_11789_),
    .ZN(_19353_));
 NOR2_X1 _36090_ (.A1(_14677_),
    .A2(_19353_),
    .ZN(_15509_));
 AND2_X1 _36091_ (.A1(_11719_),
    .A2(_11785_),
    .ZN(_15525_));
 AND2_X1 _36092_ (.A1(_11787_),
    .A2(_11788_),
    .ZN(_15524_));
 AND2_X1 _36093_ (.A1(_11786_),
    .A2(_11784_),
    .ZN(_15523_));
 CLKBUF_X3 _36094_ (.A(_11705_),
    .Z(_11790_));
 AND2_X1 _36095_ (.A1(_11790_),
    .A2(_11778_),
    .ZN(_20760_));
 AND2_X1 _36096_ (.A1(_11723_),
    .A2(_11783_),
    .ZN(_20761_));
 AND2_X1 _36097_ (.A1(_11710_),
    .A2(_11780_),
    .ZN(_15528_));
 AND2_X1 _36098_ (.A1(_11713_),
    .A2(_11779_),
    .ZN(_15529_));
 AND2_X1 _36099_ (.A1(_11790_),
    .A2(_11783_),
    .ZN(_15551_));
 BUF_X1 _36100_ (.A(_11697_),
    .Z(_11791_));
 AND2_X1 _36101_ (.A1(_11791_),
    .A2(_11784_),
    .ZN(_15550_));
 AND2_X1 _36102_ (.A1(_11723_),
    .A2(_11785_),
    .ZN(_15552_));
 AND2_X1 _36103_ (.A1(_11710_),
    .A2(_11778_),
    .ZN(_15555_));
 AND2_X1 _36104_ (.A1(_11713_),
    .A2(_11780_),
    .ZN(_15556_));
 AND2_X1 _36105_ (.A1(_11786_),
    .A2(_11788_),
    .ZN(_15563_));
 NOR2_X1 _36106_ (.A1(_15412_),
    .A2(_19353_),
    .ZN(_15562_));
 BUF_X1 _36107_ (.A(_11703_),
    .Z(_11792_));
 AND2_X1 _36108_ (.A1(_11792_),
    .A2(_11783_),
    .ZN(_15582_));
 AND2_X1 _36109_ (.A1(_11713_),
    .A2(_11778_),
    .ZN(_15583_));
 AND2_X1 _36110_ (.A1(_11790_),
    .A2(_11785_),
    .ZN(_15588_));
 AND2_X1 _36111_ (.A1(_11791_),
    .A2(_11788_),
    .ZN(_15587_));
 AND2_X1 _36112_ (.A1(_11723_),
    .A2(_11784_),
    .ZN(_15586_));
 AND2_X1 _36113_ (.A1(_11759_),
    .A2(_11753_),
    .ZN(_15595_));
 AND2_X1 _36114_ (.A1(_11741_),
    .A2(_11758_),
    .ZN(_15596_));
 AND2_X1 _36115_ (.A1(_11736_),
    .A2(_11757_),
    .ZN(_15597_));
 AND2_X1 _36116_ (.A1(_11790_),
    .A2(_11784_),
    .ZN(_15615_));
 AND2_X1 _36117_ (.A1(_11791_),
    .A2(_11789_),
    .ZN(_15614_));
 AND2_X1 _36118_ (.A1(_11723_),
    .A2(_11788_),
    .ZN(_15613_));
 AND2_X1 _36119_ (.A1(_11792_),
    .A2(_11785_),
    .ZN(_15618_));
 BUF_X2 _36120_ (.A(_11712_),
    .Z(_11793_));
 AND2_X1 _36121_ (.A1(_11793_),
    .A2(_11783_),
    .ZN(_15619_));
 AND2_X1 _36122_ (.A1(_11790_),
    .A2(_11788_),
    .ZN(_15626_));
 NOR2_X1 _36123_ (.A1(_15651_),
    .A2(_19353_),
    .ZN(_15627_));
 AND2_X1 _36124_ (.A1(_11792_),
    .A2(_11784_),
    .ZN(_15635_));
 AND2_X1 _36125_ (.A1(_11793_),
    .A2(_11785_),
    .ZN(_15634_));
 AND2_X1 _36126_ (.A1(_11793_),
    .A2(_11784_),
    .ZN(_15644_));
 AND2_X1 _36127_ (.A1(_11792_),
    .A2(_11789_),
    .ZN(_15659_));
 AND2_X1 _36128_ (.A1(_11793_),
    .A2(_11788_),
    .ZN(_15660_));
 INV_X1 _36129_ (.A(_11712_),
    .ZN(_18805_));
 NOR2_X1 _36130_ (.A1(_18805_),
    .A2(_19353_),
    .ZN(_15677_));
 BUF_X2 _36131_ (.A(net180),
    .Z(_11794_));
 AND2_X1 _36132_ (.A1(_11732_),
    .A2(_11794_),
    .ZN(_21092_));
 BUF_X2 _36133_ (.A(net179),
    .Z(_11795_));
 AND2_X1 _36134_ (.A1(_11741_),
    .A2(_11795_),
    .ZN(_21093_));
 AND2_X1 _36135_ (.A1(_11791_),
    .A2(_11717_),
    .ZN(_15687_));
 AND2_X1 _36136_ (.A1(_11694_),
    .A2(_11706_),
    .ZN(_15688_));
 CLKBUF_X3 _36137_ (.A(_11708_),
    .Z(_11796_));
 AND2_X1 _36138_ (.A1(_11796_),
    .A2(_11714_),
    .ZN(_15689_));
 AND2_X1 _36139_ (.A1(_11699_),
    .A2(_11703_),
    .ZN(_15693_));
 AND2_X1 _36140_ (.A1(_11696_),
    .A2(_11712_),
    .ZN(_15692_));
 NOR2_X1 _36141_ (.A1(_18805_),
    .A2(_19165_),
    .ZN(_15705_));
 AND2_X1 _36142_ (.A1(_11694_),
    .A2(_11703_),
    .ZN(_15754_));
 AND2_X1 _36143_ (.A1(_11699_),
    .A2(_11712_),
    .ZN(_15755_));
 NOR2_X1 _36144_ (.A1(_16722_),
    .A2(_18805_),
    .ZN(_16478_));
 CLKBUF_X3 _36145_ (.A(_11765_),
    .Z(_11797_));
 BUF_X2 _36146_ (.A(net109),
    .Z(_11798_));
 AND2_X1 _36147_ (.A1(_11797_),
    .A2(_11798_),
    .ZN(_21113_));
 BUF_X1 _36148_ (.A(net108),
    .Z(_11799_));
 AND2_X1 _36149_ (.A1(_11763_),
    .A2(_11799_),
    .ZN(_21112_));
 CLKBUF_X3 _36150_ (.A(b[19]),
    .Z(_11800_));
 AND2_X1 _36151_ (.A1(_11799_),
    .A2(_11800_),
    .ZN(_20767_));
 AND2_X1 _36152_ (.A1(_11763_),
    .A2(_11798_),
    .ZN(_20768_));
 AND2_X1 _36153_ (.A1(_11798_),
    .A2(_11800_),
    .ZN(_20770_));
 BUF_X1 _36154_ (.A(net240),
    .Z(_11801_));
 BUF_X1 _36155_ (.A(_11801_),
    .Z(_11802_));
 AND2_X1 _36156_ (.A1(_11799_),
    .A2(_11802_),
    .ZN(_20771_));
 BUF_X1 _36157_ (.A(net238),
    .Z(_11803_));
 CLKBUF_X3 _36158_ (.A(_11803_),
    .Z(_11804_));
 BUF_X2 _36159_ (.A(net113),
    .Z(_11805_));
 AND2_X1 _36160_ (.A1(_11804_),
    .A2(_11805_),
    .ZN(_15710_));
 BUF_X2 _36161_ (.A(net111),
    .Z(_11806_));
 AND2_X1 _36162_ (.A1(_11763_),
    .A2(_11806_),
    .ZN(_15709_));
 BUF_X2 _36163_ (.A(net112),
    .Z(_11807_));
 AND2_X1 _36164_ (.A1(_11797_),
    .A2(_11807_),
    .ZN(_15708_));
 AND2_X1 _36165_ (.A1(_11763_),
    .A2(_11807_),
    .ZN(_20773_));
 AND2_X1 _36166_ (.A1(_11797_),
    .A2(_11805_),
    .ZN(_20774_));
 AND2_X1 _36167_ (.A1(_11806_),
    .A2(_11800_),
    .ZN(_15713_));
 BUF_X1 _36168_ (.A(net241),
    .Z(_11808_));
 BUF_X2 _36169_ (.A(_11808_),
    .Z(_11809_));
 AND2_X1 _36170_ (.A1(_11799_),
    .A2(_11809_),
    .ZN(_15714_));
 AND2_X1 _36171_ (.A1(_11798_),
    .A2(_11802_),
    .ZN(_15715_));
 AND2_X1 _36172_ (.A1(_11763_),
    .A2(_11805_),
    .ZN(_15723_));
 AND2_X1 _36173_ (.A1(_11806_),
    .A2(_11802_),
    .ZN(_15724_));
 BUF_X2 _36174_ (.A(_11800_),
    .Z(_11810_));
 AND2_X1 _36175_ (.A1(_11810_),
    .A2(_11807_),
    .ZN(_15725_));
 AND2_X1 _36176_ (.A1(_11798_),
    .A2(_11809_),
    .ZN(_20775_));
 BUF_X4 _36177_ (.A(b[22]),
    .Z(_11811_));
 BUF_X2 _36178_ (.A(_11811_),
    .Z(_11812_));
 AND2_X1 _36179_ (.A1(_11799_),
    .A2(_11812_),
    .ZN(_20776_));
 BUF_X2 _36180_ (.A(net196),
    .Z(_11813_));
 AND2_X1 _36181_ (.A1(_11669_),
    .A2(_11813_),
    .ZN(_21095_));
 BUF_X1 _36182_ (.A(net195),
    .Z(_11814_));
 AND2_X1 _36183_ (.A1(_11664_),
    .A2(_11814_),
    .ZN(_21094_));
 BUF_X1 _36184_ (.A(_11762_),
    .Z(_11815_));
 BUF_X2 _36185_ (.A(net114),
    .Z(_11816_));
 AND2_X1 _36186_ (.A1(_11815_),
    .A2(_11816_),
    .ZN(_15736_));
 BUF_X2 _36187_ (.A(net116),
    .Z(_11817_));
 AND2_X1 _36188_ (.A1(_11804_),
    .A2(_11817_),
    .ZN(_15737_));
 BUF_X2 _36189_ (.A(net115),
    .Z(_11818_));
 AND2_X1 _36190_ (.A1(_11797_),
    .A2(_11818_),
    .ZN(_15738_));
 AND2_X1 _36191_ (.A1(_11807_),
    .A2(_11802_),
    .ZN(_20779_));
 AND2_X1 _36192_ (.A1(_11810_),
    .A2(_11805_),
    .ZN(_20778_));
 BUF_X1 _36193_ (.A(net242),
    .Z(_11819_));
 BUF_X2 _36194_ (.A(_11819_),
    .Z(_11820_));
 AND2_X1 _36195_ (.A1(_11799_),
    .A2(_11820_),
    .ZN(_15745_));
 AND2_X1 _36196_ (.A1(_11806_),
    .A2(_11809_),
    .ZN(_15746_));
 AND2_X1 _36197_ (.A1(_11798_),
    .A2(_11812_),
    .ZN(_15747_));
 AND2_X1 _36198_ (.A1(_11790_),
    .A2(_11714_),
    .ZN(_15763_));
 NOR2_X1 _36199_ (.A1(_15651_),
    .A2(_19165_),
    .ZN(_15764_));
 AND2_X1 _36200_ (.A1(_11806_),
    .A2(_11812_),
    .ZN(_15780_));
 BUF_X1 _36201_ (.A(net243),
    .Z(_11821_));
 BUF_X1 _36202_ (.A(_11821_),
    .Z(_11822_));
 AND2_X1 _36203_ (.A1(_11799_),
    .A2(_11822_),
    .ZN(_15781_));
 AND2_X1 _36204_ (.A1(_11798_),
    .A2(_11820_),
    .ZN(_15782_));
 AND2_X1 _36205_ (.A1(_11797_),
    .A2(_11817_),
    .ZN(_20781_));
 AND2_X1 _36206_ (.A1(_11815_),
    .A2(_11818_),
    .ZN(_20782_));
 AND2_X1 _36207_ (.A1(_11807_),
    .A2(_11809_),
    .ZN(_15787_));
 AND2_X1 _36208_ (.A1(_11810_),
    .A2(_11816_),
    .ZN(_15786_));
 BUF_X2 _36209_ (.A(_11801_),
    .Z(_11823_));
 AND2_X1 _36210_ (.A1(_11823_),
    .A2(_11805_),
    .ZN(_15785_));
 AND2_X1 _36211_ (.A1(_11806_),
    .A2(_11820_),
    .ZN(_15801_));
 AND2_X1 _36212_ (.A1(_11805_),
    .A2(_11809_),
    .ZN(_15803_));
 AND2_X1 _36213_ (.A1(_11807_),
    .A2(_11811_),
    .ZN(_15802_));
 AND2_X1 _36214_ (.A1(_11798_),
    .A2(_11822_),
    .ZN(_20785_));
 BUF_X1 _36215_ (.A(b[25]),
    .Z(_11824_));
 BUF_X2 _36216_ (.A(_11824_),
    .Z(_11825_));
 AND2_X1 _36217_ (.A1(_11799_),
    .A2(_11825_),
    .ZN(_20784_));
 AND2_X1 _36218_ (.A1(_11815_),
    .A2(_11817_),
    .ZN(_15811_));
 AND2_X1 _36219_ (.A1(_11823_),
    .A2(_11816_),
    .ZN(_15812_));
 AND2_X1 _36220_ (.A1(_11810_),
    .A2(_11818_),
    .ZN(_15813_));
 AND2_X1 _36221_ (.A1(_11805_),
    .A2(_11811_),
    .ZN(_20787_));
 AND2_X1 _36222_ (.A1(_11807_),
    .A2(_11820_),
    .ZN(_20788_));
 AND2_X1 _36223_ (.A1(_11806_),
    .A2(_11822_),
    .ZN(_15827_));
 AND2_X1 _36224_ (.A1(_11798_),
    .A2(_11825_),
    .ZN(_15828_));
 AND2_X1 _36225_ (.A1(_11810_),
    .A2(_11817_),
    .ZN(_15835_));
 AND2_X1 _36226_ (.A1(_11816_),
    .A2(_11809_),
    .ZN(_15836_));
 AND2_X1 _36227_ (.A1(_11823_),
    .A2(_11818_),
    .ZN(_15837_));
 BUF_X2 _36228_ (.A(net117),
    .Z(_11826_));
 AND2_X1 _36229_ (.A1(_11815_),
    .A2(_11826_),
    .ZN(_15840_));
 INV_X4 _36230_ (.A(_11765_),
    .ZN(_15870_));
 BUF_X2 _36231_ (.A(a[217]),
    .Z(_11827_));
 INV_X2 _36232_ (.A(_11827_),
    .ZN(_19303_));
 NOR2_X1 _36233_ (.A1(_15870_),
    .A2(_19303_),
    .ZN(_15841_));
 BUF_X2 _36234_ (.A(_11808_),
    .Z(_11828_));
 AND2_X1 _36235_ (.A1(_11828_),
    .A2(_11818_),
    .ZN(_15857_));
 AND2_X1 _36236_ (.A1(_11810_),
    .A2(_11826_),
    .ZN(_15858_));
 AND2_X1 _36237_ (.A1(_11823_),
    .A2(_11817_),
    .ZN(_15856_));
 AND2_X1 _36238_ (.A1(_11816_),
    .A2(_11811_),
    .ZN(_20791_));
 AND2_X1 _36239_ (.A1(_11805_),
    .A2(_11820_),
    .ZN(_20790_));
 AND2_X1 _36240_ (.A1(_11807_),
    .A2(_11822_),
    .ZN(_15861_));
 AND2_X1 _36241_ (.A1(_11806_),
    .A2(_11825_),
    .ZN(_15862_));
 AND2_X1 _36242_ (.A1(_11805_),
    .A2(_11821_),
    .ZN(_15884_));
 AND2_X1 _36243_ (.A1(_11807_),
    .A2(_11825_),
    .ZN(_15883_));
 AND2_X1 _36244_ (.A1(_11828_),
    .A2(_11817_),
    .ZN(_15892_));
 AND2_X1 _36245_ (.A1(_11816_),
    .A2(_11820_),
    .ZN(_15891_));
 BUF_X2 _36246_ (.A(_11811_),
    .Z(_11829_));
 AND2_X1 _36247_ (.A1(_11829_),
    .A2(_11818_),
    .ZN(_15890_));
 AND2_X1 _36248_ (.A1(_11823_),
    .A2(_11826_),
    .ZN(_15895_));
 INV_X4 _36249_ (.A(_11800_),
    .ZN(_15915_));
 NOR2_X1 _36250_ (.A1(_15915_),
    .A2(_19303_),
    .ZN(_15896_));
 AND2_X1 _36251_ (.A1(_11816_),
    .A2(_11821_),
    .ZN(_15911_));
 AND2_X1 _36252_ (.A1(_11805_),
    .A2(_11825_),
    .ZN(_15912_));
 AND2_X1 _36253_ (.A1(_11818_),
    .A2(_11820_),
    .ZN(_15921_));
 AND2_X1 _36254_ (.A1(_11828_),
    .A2(_11826_),
    .ZN(_15920_));
 AND2_X1 _36255_ (.A1(_11829_),
    .A2(_11817_),
    .ZN(_15922_));
 AND2_X1 _36256_ (.A1(_11828_),
    .A2(_11827_),
    .ZN(_15931_));
 AND2_X1 _36257_ (.A1(_11817_),
    .A2(_11820_),
    .ZN(_15930_));
 AND2_X1 _36258_ (.A1(_11829_),
    .A2(_11826_),
    .ZN(_15929_));
 AND2_X1 _36259_ (.A1(_11818_),
    .A2(_11821_),
    .ZN(_15934_));
 AND2_X1 _36260_ (.A1(_11816_),
    .A2(_11825_),
    .ZN(_15935_));
 AND2_X1 _36261_ (.A1(_11817_),
    .A2(_11821_),
    .ZN(_15947_));
 AND2_X1 _36262_ (.A1(_11818_),
    .A2(_11824_),
    .ZN(_15948_));
 CLKBUF_X3 _36263_ (.A(_11819_),
    .Z(_11830_));
 AND2_X1 _36264_ (.A1(_11830_),
    .A2(_11826_),
    .ZN(_15956_));
 INV_X4 _36265_ (.A(_11811_),
    .ZN(_15964_));
 NOR2_X1 _36266_ (.A1(_15964_),
    .A2(_19303_),
    .ZN(_15957_));
 AND2_X1 _36267_ (.A1(_11817_),
    .A2(_11824_),
    .ZN(_15969_));
 BUF_X1 _36268_ (.A(_11821_),
    .Z(_11831_));
 AND2_X1 _36269_ (.A1(_11831_),
    .A2(_11827_),
    .ZN(_15980_));
 AND2_X1 _36270_ (.A1(_11826_),
    .A2(_11824_),
    .ZN(_15981_));
 INV_X1 _36271_ (.A(_11824_),
    .ZN(_18757_));
 NOR2_X1 _36272_ (.A1(_18757_),
    .A2(_19303_),
    .ZN(_15984_));
 BUF_X2 _36273_ (.A(net53),
    .Z(_11832_));
 AND2_X1 _36274_ (.A1(_11830_),
    .A2(_11832_),
    .ZN(_15987_));
 BUF_X2 _36275_ (.A(a[153]),
    .Z(_11833_));
 INV_X2 _36276_ (.A(_11833_),
    .ZN(_19122_));
 NOR2_X1 _36277_ (.A1(_15964_),
    .A2(_19122_),
    .ZN(_15988_));
 BUF_X2 _36278_ (.A(net51),
    .Z(_11834_));
 AND2_X1 _36279_ (.A1(_11830_),
    .A2(_11834_),
    .ZN(_16029_));
 AND2_X1 _36280_ (.A1(_11828_),
    .A2(_11832_),
    .ZN(_16030_));
 BUF_X2 _36281_ (.A(net52),
    .Z(_11835_));
 AND2_X1 _36282_ (.A1(_11829_),
    .A2(_11835_),
    .ZN(_16031_));
 BUF_X2 _36283_ (.A(net49),
    .Z(_11836_));
 AND2_X1 _36284_ (.A1(_11831_),
    .A2(_11836_),
    .ZN(_16022_));
 CLKBUF_X3 _36285_ (.A(_11824_),
    .Z(_11837_));
 BUF_X2 _36286_ (.A(net48),
    .Z(_11838_));
 AND2_X1 _36287_ (.A1(_11837_),
    .A2(_11838_),
    .ZN(_16023_));
 AND2_X1 _36288_ (.A1(_11831_),
    .A2(_11838_),
    .ZN(_16019_));
 BUF_X2 _36289_ (.A(net47),
    .Z(_11839_));
 AND2_X1 _36290_ (.A1(_11837_),
    .A2(_11839_),
    .ZN(_16018_));
 AND2_X1 _36291_ (.A1(_11828_),
    .A2(_11833_),
    .ZN(_15993_));
 AND2_X1 _36292_ (.A1(_11830_),
    .A2(_11835_),
    .ZN(_15992_));
 AND2_X1 _36293_ (.A1(_11829_),
    .A2(_11832_),
    .ZN(_15991_));
 AND2_X1 _36294_ (.A1(_11831_),
    .A2(_11834_),
    .ZN(_15996_));
 AND2_X1 _36295_ (.A1(_11837_),
    .A2(_11836_),
    .ZN(_15997_));
 AND2_X1 _36296_ (.A1(_11831_),
    .A2(_11835_),
    .ZN(_16006_));
 AND2_X1 _36297_ (.A1(_11837_),
    .A2(_11834_),
    .ZN(_16005_));
 AND2_X1 _36298_ (.A1(_11828_),
    .A2(_11835_),
    .ZN(_16054_));
 AND2_X1 _36299_ (.A1(_11830_),
    .A2(_11836_),
    .ZN(_16053_));
 AND2_X1 _36300_ (.A1(_11829_),
    .A2(_11834_),
    .ZN(_16052_));
 AND2_X1 _36301_ (.A1(_11831_),
    .A2(_11839_),
    .ZN(_16041_));
 BUF_X2 _36302_ (.A(net46),
    .Z(_11840_));
 AND2_X1 _36303_ (.A1(_11837_),
    .A2(_11840_),
    .ZN(_16042_));
 AND2_X1 _36304_ (.A1(_11830_),
    .A2(_11838_),
    .ZN(_20795_));
 AND2_X1 _36305_ (.A1(_11829_),
    .A2(_11836_),
    .ZN(_20794_));
 AND2_X1 _36306_ (.A1(_11823_),
    .A2(_11832_),
    .ZN(_16057_));
 NOR2_X1 _36307_ (.A1(_15915_),
    .A2(_19122_),
    .ZN(_16058_));
 BUF_X2 _36308_ (.A(_11819_),
    .Z(_11841_));
 AND2_X1 _36309_ (.A1(_11841_),
    .A2(_11839_),
    .ZN(_20797_));
 AND2_X1 _36310_ (.A1(_11829_),
    .A2(_11838_),
    .ZN(_20796_));
 AND2_X1 _36311_ (.A1(_11810_),
    .A2(_11832_),
    .ZN(_16080_));
 AND2_X1 _36312_ (.A1(_11828_),
    .A2(_11834_),
    .ZN(_16081_));
 BUF_X1 _36313_ (.A(_11801_),
    .Z(_11842_));
 AND2_X1 _36314_ (.A1(_11842_),
    .A2(_11835_),
    .ZN(_16082_));
 AND2_X1 _36315_ (.A1(_11831_),
    .A2(_11840_),
    .ZN(_16072_));
 BUF_X2 _36316_ (.A(net45),
    .Z(_11843_));
 AND2_X1 _36317_ (.A1(_11837_),
    .A2(_11843_),
    .ZN(_16073_));
 AND2_X1 _36318_ (.A1(_11831_),
    .A2(_11843_),
    .ZN(_20801_));
 AND2_X1 _36319_ (.A1(_11810_),
    .A2(_11835_),
    .ZN(_16106_));
 AND2_X1 _36320_ (.A1(_11828_),
    .A2(_11836_),
    .ZN(_16105_));
 AND2_X1 _36321_ (.A1(_11842_),
    .A2(_11834_),
    .ZN(_16104_));
 AND2_X1 _36322_ (.A1(_11815_),
    .A2(_11832_),
    .ZN(_16109_));
 NOR2_X1 _36323_ (.A1(_15870_),
    .A2(_19122_),
    .ZN(_16110_));
 AND2_X1 _36324_ (.A1(_11828_),
    .A2(_11838_),
    .ZN(_16124_));
 AND2_X1 _36325_ (.A1(_11841_),
    .A2(_11840_),
    .ZN(_16125_));
 AND2_X1 _36326_ (.A1(_11829_),
    .A2(_11839_),
    .ZN(_16126_));
 AND2_X1 _36327_ (.A1(_11842_),
    .A2(_11836_),
    .ZN(_16133_));
 AND2_X1 _36328_ (.A1(_11815_),
    .A2(_11835_),
    .ZN(_16134_));
 AND2_X1 _36329_ (.A1(_11810_),
    .A2(_11834_),
    .ZN(_16135_));
 BUF_X1 _36330_ (.A(net44),
    .Z(_11844_));
 AND2_X1 _36331_ (.A1(_11831_),
    .A2(_11844_),
    .ZN(_16151_));
 AND2_X1 _36332_ (.A1(_11829_),
    .A2(_11840_),
    .ZN(_16150_));
 AND2_X1 _36333_ (.A1(_11841_),
    .A2(_11843_),
    .ZN(_16152_));
 AND2_X1 _36334_ (.A1(_11815_),
    .A2(_11834_),
    .ZN(_20804_));
 AND2_X1 _36335_ (.A1(_11797_),
    .A2(_11835_),
    .ZN(_20805_));
 BUF_X2 _36336_ (.A(_11808_),
    .Z(_11845_));
 AND2_X1 _36337_ (.A1(_11845_),
    .A2(_11839_),
    .ZN(_16156_));
 AND2_X1 _36338_ (.A1(_11810_),
    .A2(_11836_),
    .ZN(_16155_));
 AND2_X1 _36339_ (.A1(_11842_),
    .A2(_11838_),
    .ZN(_16154_));
 BUF_X2 _36340_ (.A(net213),
    .Z(_11846_));
 AND2_X1 _36341_ (.A1(_11797_),
    .A2(_11846_),
    .ZN(_21096_));
 BUF_X1 _36342_ (.A(net212),
    .Z(_11847_));
 AND2_X1 _36343_ (.A1(_11815_),
    .A2(_11847_),
    .ZN(_21097_));
 AND2_X1 _36344_ (.A1(_11842_),
    .A2(_11839_),
    .ZN(_20807_));
 BUF_X2 _36345_ (.A(_11800_),
    .Z(_11848_));
 AND2_X1 _36346_ (.A1(_11848_),
    .A2(_11838_),
    .ZN(_20808_));
 AND2_X1 _36347_ (.A1(_11845_),
    .A2(_11840_),
    .ZN(_16171_));
 AND2_X1 _36348_ (.A1(_11841_),
    .A2(_11844_),
    .ZN(_16170_));
 BUF_X2 _36349_ (.A(_11811_),
    .Z(_11849_));
 AND2_X1 _36350_ (.A1(_11849_),
    .A2(_11843_),
    .ZN(_16172_));
 AND2_X1 _36351_ (.A1(_11804_),
    .A2(_11835_),
    .ZN(_16185_));
 AND2_X1 _36352_ (.A1(_11815_),
    .A2(_11836_),
    .ZN(_16184_));
 AND2_X1 _36353_ (.A1(_11797_),
    .A2(_11834_),
    .ZN(_16183_));
 AND2_X1 _36354_ (.A1(_11845_),
    .A2(_11843_),
    .ZN(_20809_));
 AND2_X1 _36355_ (.A1(_11849_),
    .A2(_11844_),
    .ZN(_20810_));
 AND2_X1 _36356_ (.A1(_11815_),
    .A2(_11838_),
    .ZN(_16197_));
 AND2_X1 _36357_ (.A1(_11842_),
    .A2(_11840_),
    .ZN(_16198_));
 AND2_X1 _36358_ (.A1(_11848_),
    .A2(_11839_),
    .ZN(_16199_));
 AND2_X1 _36359_ (.A1(_11845_),
    .A2(_11844_),
    .ZN(_16212_));
 AND2_X1 _36360_ (.A1(_11848_),
    .A2(_11840_),
    .ZN(_16211_));
 AND2_X1 _36361_ (.A1(_11842_),
    .A2(_11843_),
    .ZN(_16210_));
 AND2_X1 _36362_ (.A1(_11797_),
    .A2(_11838_),
    .ZN(_20813_));
 BUF_X1 _36363_ (.A(_11762_),
    .Z(_11850_));
 AND2_X1 _36364_ (.A1(_11850_),
    .A2(_11839_),
    .ZN(_20814_));
 AND2_X1 _36365_ (.A1(_11848_),
    .A2(_11843_),
    .ZN(_20816_));
 AND2_X1 _36366_ (.A1(_11842_),
    .A2(_11844_),
    .ZN(_20817_));
 BUF_X1 _36367_ (.A(_11803_),
    .Z(_11851_));
 AND2_X1 _36368_ (.A1(_11851_),
    .A2(_11838_),
    .ZN(_16221_));
 AND2_X1 _36369_ (.A1(_11850_),
    .A2(_11840_),
    .ZN(_16220_));
 AND2_X1 _36370_ (.A1(_11797_),
    .A2(_11839_),
    .ZN(_16219_));
 AND2_X1 _36371_ (.A1(_11848_),
    .A2(_11844_),
    .ZN(_20818_));
 AND2_X1 _36372_ (.A1(_11850_),
    .A2(_11843_),
    .ZN(_20819_));
 CLKBUF_X3 _36373_ (.A(_11765_),
    .Z(_11852_));
 AND2_X1 _36374_ (.A1(_11852_),
    .A2(_11840_),
    .ZN(_19127_));
 AND2_X1 _36375_ (.A1(_11851_),
    .A2(_11839_),
    .ZN(_19126_));
 AND2_X1 _36376_ (.A1(_11850_),
    .A2(_11844_),
    .ZN(_21105_));
 AND2_X1 _36377_ (.A1(_11852_),
    .A2(_11843_),
    .ZN(_21104_));
 BUF_X2 _36378_ (.A(_11662_),
    .Z(_11853_));
 BUF_X1 _36379_ (.A(net92),
    .Z(_11854_));
 AND2_X1 _36380_ (.A1(_11853_),
    .A2(_11854_),
    .ZN(_20820_));
 BUF_X2 _36381_ (.A(net93),
    .Z(_11855_));
 AND2_X1 _36382_ (.A1(_11664_),
    .A2(_11855_),
    .ZN(_20821_));
 AND2_X1 _36383_ (.A1(_11853_),
    .A2(_11855_),
    .ZN(_20823_));
 AND2_X1 _36384_ (.A1(_11747_),
    .A2(_11854_),
    .ZN(_20824_));
 BUF_X2 _36385_ (.A(net94),
    .Z(_11856_));
 AND2_X1 _36386_ (.A1(_11664_),
    .A2(_11856_),
    .ZN(_16226_));
 BUF_X1 _36387_ (.A(_11667_),
    .Z(_11857_));
 BUF_X2 _36388_ (.A(net96),
    .Z(_11858_));
 AND2_X1 _36389_ (.A1(_11857_),
    .A2(_11858_),
    .ZN(_16225_));
 BUF_X2 _36390_ (.A(net95),
    .Z(_11859_));
 AND2_X1 _36391_ (.A1(_11669_),
    .A2(_11859_),
    .ZN(_16224_));
 BUF_X1 _36392_ (.A(_11656_),
    .Z(_11860_));
 AND2_X1 _36393_ (.A1(_11860_),
    .A2(_11859_),
    .ZN(_20826_));
 AND2_X1 _36394_ (.A1(_11669_),
    .A2(_11858_),
    .ZN(_20827_));
 AND2_X1 _36395_ (.A1(_11853_),
    .A2(_11856_),
    .ZN(_16231_));
 AND2_X1 _36396_ (.A1(_11666_),
    .A2(_11854_),
    .ZN(_16230_));
 AND2_X1 _36397_ (.A1(_11747_),
    .A2(_11855_),
    .ZN(_16229_));
 AND2_X1 _36398_ (.A1(_11769_),
    .A2(_11854_),
    .ZN(_20828_));
 AND2_X1 _36399_ (.A1(_11666_),
    .A2(_11855_),
    .ZN(_20829_));
 AND2_X1 _36400_ (.A1(_11747_),
    .A2(_11856_),
    .ZN(_16244_));
 AND2_X1 _36401_ (.A1(_11860_),
    .A2(_11858_),
    .ZN(_16245_));
 AND2_X1 _36402_ (.A1(_11853_),
    .A2(_11859_),
    .ZN(_16246_));
 AND2_X1 _36403_ (.A1(_11747_),
    .A2(_11859_),
    .ZN(_20831_));
 AND2_X1 _36404_ (.A1(_11853_),
    .A2(_11858_),
    .ZN(_20832_));
 AND2_X1 _36405_ (.A1(_11748_),
    .A2(_11854_),
    .ZN(_16252_));
 AND2_X1 _36406_ (.A1(_11666_),
    .A2(_11856_),
    .ZN(_16253_));
 AND2_X1 _36407_ (.A1(_11769_),
    .A2(_11855_),
    .ZN(_16254_));
 BUF_X2 _36408_ (.A(net97),
    .Z(_11861_));
 AND2_X1 _36409_ (.A1(_11860_),
    .A2(_11861_),
    .ZN(_16261_));
 BUF_X2 _36410_ (.A(a[199]),
    .Z(_11862_));
 AND2_X1 _36411_ (.A1(_11857_),
    .A2(_11862_),
    .ZN(_16262_));
 BUF_X2 _36412_ (.A(net98),
    .Z(_11863_));
 AND2_X1 _36413_ (.A1(_11669_),
    .A2(_11863_),
    .ZN(_16263_));
 INV_X2 _36414_ (.A(_11862_),
    .ZN(_16485_));
 NOR2_X1 _36415_ (.A1(_15313_),
    .A2(_16485_),
    .ZN(_20834_));
 AND2_X1 _36416_ (.A1(_11860_),
    .A2(_11863_),
    .ZN(_20835_));
 AND2_X1 _36417_ (.A1(_11769_),
    .A2(_11856_),
    .ZN(_16270_));
 AND2_X1 _36418_ (.A1(_11749_),
    .A2(_11854_),
    .ZN(_16271_));
 AND2_X1 _36419_ (.A1(_11748_),
    .A2(_11855_),
    .ZN(_16272_));
 AND2_X1 _36420_ (.A1(_11853_),
    .A2(_11861_),
    .ZN(_16277_));
 AND2_X1 _36421_ (.A1(_11666_),
    .A2(_11859_),
    .ZN(_16276_));
 AND2_X1 _36422_ (.A1(_11747_),
    .A2(_11858_),
    .ZN(_16275_));
 AND2_X1 _36423_ (.A1(_11702_),
    .A2(_11716_),
    .ZN(_20838_));
 AND2_X1 _36424_ (.A1(_11787_),
    .A2(_11722_),
    .ZN(_20839_));
 AND2_X1 _36425_ (.A1(_11749_),
    .A2(_11855_),
    .ZN(_20842_));
 AND2_X1 _36426_ (.A1(_11750_),
    .A2(_11854_),
    .ZN(_20841_));
 BUF_X2 _36427_ (.A(_11650_),
    .Z(_11864_));
 AND2_X1 _36428_ (.A1(_11864_),
    .A2(_11856_),
    .ZN(_16299_));
 AND2_X1 _36429_ (.A1(_11666_),
    .A2(_11858_),
    .ZN(_16300_));
 AND2_X1 _36430_ (.A1(_11769_),
    .A2(_11859_),
    .ZN(_16301_));
 AND2_X1 _36431_ (.A1(_11860_),
    .A2(_11862_),
    .ZN(_16306_));
 BUF_X2 _36432_ (.A(_11659_),
    .Z(_11865_));
 AND2_X1 _36433_ (.A1(_11865_),
    .A2(_11861_),
    .ZN(_16305_));
 AND2_X1 _36434_ (.A1(_11853_),
    .A2(_11863_),
    .ZN(_16304_));
 NOR2_X1 _36435_ (.A1(_15238_),
    .A2(_16485_),
    .ZN(_16322_));
 BUF_X2 _36436_ (.A(_11647_),
    .Z(_11866_));
 AND2_X1 _36437_ (.A1(_11866_),
    .A2(_11861_),
    .ZN(_16321_));
 AND2_X1 _36438_ (.A1(_11865_),
    .A2(_11863_),
    .ZN(_16320_));
 AND2_X1 _36439_ (.A1(_11769_),
    .A2(_11858_),
    .ZN(_20844_));
 AND2_X1 _36440_ (.A1(_11864_),
    .A2(_11859_),
    .ZN(_20845_));
 BUF_X1 _36441_ (.A(_11645_),
    .Z(_11867_));
 AND2_X1 _36442_ (.A1(_11867_),
    .A2(_11856_),
    .ZN(_16325_));
 AND2_X1 _36443_ (.A1(_11750_),
    .A2(_11855_),
    .ZN(_16326_));
 BUF_X2 _36444_ (.A(net101),
    .Z(_11868_));
 AND2_X1 _36445_ (.A1(_11860_),
    .A2(_11868_),
    .ZN(_16334_));
 BUF_X2 _36446_ (.A(a[201]),
    .Z(_11869_));
 INV_X2 _36447_ (.A(_11869_),
    .ZN(_19253_));
 NOR2_X1 _36448_ (.A1(_15313_),
    .A2(_19253_),
    .ZN(_16333_));
 AND2_X1 _36449_ (.A1(_11853_),
    .A2(_11868_),
    .ZN(_16350_));
 AND2_X1 _36450_ (.A1(_11866_),
    .A2(_11863_),
    .ZN(_16349_));
 AND2_X1 _36451_ (.A1(_11865_),
    .A2(_11862_),
    .ZN(_16348_));
 AND2_X1 _36452_ (.A1(_11769_),
    .A2(_11861_),
    .ZN(_20847_));
 AND2_X1 _36453_ (.A1(_11864_),
    .A2(_11858_),
    .ZN(_20848_));
 AND2_X1 _36454_ (.A1(_11867_),
    .A2(_11859_),
    .ZN(_16353_));
 BUF_X2 _36455_ (.A(_11643_),
    .Z(_11870_));
 AND2_X1 _36456_ (.A1(_11870_),
    .A2(_11856_),
    .ZN(_16354_));
 AND2_X1 _36457_ (.A1(_11864_),
    .A2(_11861_),
    .ZN(_16376_));
 AND2_X1 _36458_ (.A1(_11866_),
    .A2(_11862_),
    .ZN(_16377_));
 AND2_X1 _36459_ (.A1(_11769_),
    .A2(_11863_),
    .ZN(_16378_));
 AND2_X1 _36460_ (.A1(_11867_),
    .A2(_11858_),
    .ZN(_16382_));
 AND2_X1 _36461_ (.A1(_11870_),
    .A2(_11859_),
    .ZN(_16381_));
 AND2_X1 _36462_ (.A1(_11865_),
    .A2(_11868_),
    .ZN(_16388_));
 NOR2_X1 _36463_ (.A1(_15238_),
    .A2(_19253_),
    .ZN(_16389_));
 AND2_X1 _36464_ (.A1(_11867_),
    .A2(_11861_),
    .ZN(_16413_));
 AND2_X1 _36465_ (.A1(_11870_),
    .A2(_11858_),
    .ZN(_16414_));
 AND2_X1 _36466_ (.A1(_11864_),
    .A2(_11863_),
    .ZN(_16417_));
 AND2_X1 _36467_ (.A1(_11866_),
    .A2(_11868_),
    .ZN(_16418_));
 NOR2_X1 _36468_ (.A1(_15196_),
    .A2(_16485_),
    .ZN(_16419_));
 BUF_X2 _36469_ (.A(net229),
    .Z(_11871_));
 AND2_X1 _36470_ (.A1(_11772_),
    .A2(_11871_),
    .ZN(_21099_));
 BUF_X2 _36471_ (.A(net228),
    .Z(_11872_));
 AND2_X1 _36472_ (.A1(_11782_),
    .A2(_11872_),
    .ZN(_21098_));
 AND2_X1 _36473_ (.A1(_11866_),
    .A2(_11869_),
    .ZN(_16431_));
 AND2_X1 _36474_ (.A1(_11864_),
    .A2(_11862_),
    .ZN(_16432_));
 AND2_X1 _36475_ (.A1(_11769_),
    .A2(_11868_),
    .ZN(_16433_));
 AND2_X1 _36476_ (.A1(_11867_),
    .A2(_11863_),
    .ZN(_16437_));
 AND2_X1 _36477_ (.A1(_11870_),
    .A2(_11861_),
    .ZN(_16436_));
 AND2_X1 _36478_ (.A1(_11864_),
    .A2(_11868_),
    .ZN(_16445_));
 NOR2_X1 _36479_ (.A1(_15196_),
    .A2(_19253_),
    .ZN(_16444_));
 AND2_X1 _36480_ (.A1(_11867_),
    .A2(_11862_),
    .ZN(_16452_));
 AND2_X1 _36481_ (.A1(_11870_),
    .A2(_11863_),
    .ZN(_16453_));
 NOR2_X1 _36482_ (.A1(_18713_),
    .A2(_16485_),
    .ZN(_16466_));
 NOR2_X1 _36483_ (.A1(_18713_),
    .A2(_19253_),
    .ZN(_16493_));
 BUF_X1 _36484_ (.A(_11718_),
    .Z(_11873_));
 AND2_X1 _36485_ (.A1(_11702_),
    .A2(_11873_),
    .ZN(_21106_));
 AND2_X1 _36486_ (.A1(_11722_),
    .A2(_11716_),
    .ZN(_21107_));
 NOR2_X1 _36487_ (.A1(_18757_),
    .A2(_19122_),
    .ZN(_16496_));
 BUF_X1 _36488_ (.A(_11821_),
    .Z(_11874_));
 AND2_X1 _36489_ (.A1(_11874_),
    .A2(_11833_),
    .ZN(_16504_));
 AND2_X1 _36490_ (.A1(_11837_),
    .A2(_11832_),
    .ZN(_16503_));
 AND2_X1 _36491_ (.A1(_11837_),
    .A2(_11835_),
    .ZN(_16507_));
 AND2_X1 _36492_ (.A1(_11707_),
    .A2(_11716_),
    .ZN(_16540_));
 AND2_X1 _36493_ (.A1(_11786_),
    .A2(_11711_),
    .ZN(_16539_));
 AND2_X1 _36494_ (.A1(_11787_),
    .A2(_11704_),
    .ZN(_16538_));
 BUF_X1 _36495_ (.A(_11776_),
    .Z(_11875_));
 AND2_X1 _36496_ (.A1(_11694_),
    .A2(_11875_),
    .ZN(_16518_));
 AND2_X1 _36497_ (.A1(_11696_),
    .A2(_11716_),
    .ZN(_16519_));
 AND2_X1 _36498_ (.A1(_11699_),
    .A2(_11718_),
    .ZN(_16520_));
 AND2_X1 _36499_ (.A1(_11722_),
    .A2(_11708_),
    .ZN(_20852_));
 AND2_X1 _36500_ (.A1(_11787_),
    .A2(_11707_),
    .ZN(_20856_));
 AND2_X1 _36501_ (.A1(_11786_),
    .A2(_11704_),
    .ZN(_20857_));
 AND2_X1 _36502_ (.A1(_11791_),
    .A2(_11711_),
    .ZN(_16530_));
 AND2_X1 _36503_ (.A1(_11722_),
    .A2(_11706_),
    .ZN(_16529_));
 AND2_X1 _36504_ (.A1(_11702_),
    .A2(_11708_),
    .ZN(_16528_));
 AND2_X1 _36505_ (.A1(_11787_),
    .A2(_11711_),
    .ZN(_16551_));
 AND2_X1 _36506_ (.A1(_11791_),
    .A2(_11722_),
    .ZN(_16552_));
 AND2_X1 _36507_ (.A1(_11786_),
    .A2(_11702_),
    .ZN(_16553_));
 AND2_X1 _36508_ (.A1(_11707_),
    .A2(_11718_),
    .ZN(_20862_));
 AND2_X1 _36509_ (.A1(_11704_),
    .A2(_11716_),
    .ZN(_20861_));
 BUF_X2 _36510_ (.A(net13),
    .Z(_11876_));
 AND2_X1 _36511_ (.A1(_11741_),
    .A2(_11876_),
    .ZN(_21100_));
 BUF_X2 _36512_ (.A(net14),
    .Z(_11877_));
 AND2_X1 _36513_ (.A1(_11732_),
    .A2(_11877_),
    .ZN(_21101_));
 AND2_X1 _36514_ (.A1(_11787_),
    .A2(_11702_),
    .ZN(_20864_));
 AND2_X1 _36515_ (.A1(_11786_),
    .A2(_11722_),
    .ZN(_20865_));
 AND2_X1 _36516_ (.A1(_11707_),
    .A2(_11875_),
    .ZN(_16562_));
 AND2_X1 _36517_ (.A1(_11711_),
    .A2(_11716_),
    .ZN(_16561_));
 AND2_X1 _36518_ (.A1(_11704_),
    .A2(_11718_),
    .ZN(_16560_));
 AND2_X1 _36519_ (.A1(_11860_),
    .A2(_11854_),
    .ZN(_21110_));
 AND2_X1 _36520_ (.A1(_11669_),
    .A2(_11855_),
    .ZN(_21111_));
 BUF_X2 _36521_ (.A(a[9]),
    .Z(_11878_));
 INV_X2 _36522_ (.A(_11878_),
    .ZN(_18712_));
 NOR2_X1 _36523_ (.A1(_18713_),
    .A2(_18712_),
    .ZN(_16565_));
 AND2_X1 _36524_ (.A1(_11867_),
    .A2(_11878_),
    .ZN(_18638_));
 BUF_X2 _36525_ (.A(net221),
    .Z(_11879_));
 AND2_X1 _36526_ (.A1(_11870_),
    .A2(_11879_),
    .ZN(_18637_));
 BUF_X2 _36527_ (.A(net211),
    .Z(_11880_));
 AND2_X1 _36528_ (.A1(_11867_),
    .A2(_11880_),
    .ZN(_17644_));
 BUF_X2 _36529_ (.A(net201),
    .Z(_11881_));
 AND2_X1 _36530_ (.A1(_11870_),
    .A2(_11881_),
    .ZN(_17645_));
 AND2_X1 _36531_ (.A1(_11870_),
    .A2(_11880_),
    .ZN(_17641_));
 BUF_X2 _36532_ (.A(net181),
    .Z(_11882_));
 AND2_X1 _36533_ (.A1(_11867_),
    .A2(_11882_),
    .ZN(_16569_));
 BUF_X2 _36534_ (.A(net171),
    .Z(_11883_));
 AND2_X1 _36535_ (.A1(_11870_),
    .A2(_11883_),
    .ZN(_16568_));
 AND2_X1 _36536_ (.A1(_11867_),
    .A2(_11883_),
    .ZN(_16577_));
 BUF_X2 _36537_ (.A(net160),
    .Z(_11884_));
 AND2_X1 _36538_ (.A1(_11870_),
    .A2(_11884_),
    .ZN(_16578_));
 AND2_X1 _36539_ (.A1(_11864_),
    .A2(_11882_),
    .ZN(_20867_));
 BUF_X2 _36540_ (.A(_11653_),
    .Z(_11885_));
 BUF_X2 _36541_ (.A(net190),
    .Z(_11886_));
 AND2_X1 _36542_ (.A1(_11885_),
    .A2(_11886_),
    .ZN(_20868_));
 AND2_X1 _36543_ (.A1(_11864_),
    .A2(_11886_),
    .ZN(_16583_));
 AND2_X1 _36544_ (.A1(_11866_),
    .A2(_11880_),
    .ZN(_16582_));
 AND2_X1 _36545_ (.A1(_11885_),
    .A2(_11881_),
    .ZN(_16581_));
 AND2_X1 _36546_ (.A1(_11865_),
    .A2(_11879_),
    .ZN(_16589_));
 NOR2_X1 _36547_ (.A1(_15238_),
    .A2(_18712_),
    .ZN(_16590_));
 AND2_X1 _36548_ (.A1(_11853_),
    .A2(_11879_),
    .ZN(_16624_));
 AND2_X1 _36549_ (.A1(_11866_),
    .A2(_11881_),
    .ZN(_16623_));
 AND2_X1 _36550_ (.A1(_11865_),
    .A2(_11880_),
    .ZN(_16622_));
 AND2_X1 _36551_ (.A1(_11864_),
    .A2(_11883_),
    .ZN(_20872_));
 BUF_X1 _36552_ (.A(_11645_),
    .Z(_11887_));
 AND2_X1 _36553_ (.A1(_11887_),
    .A2(_11884_),
    .ZN(_16618_));
 BUF_X2 _36554_ (.A(_11643_),
    .Z(_11888_));
 AND2_X1 _36555_ (.A1(_11888_),
    .A2(_11686_),
    .ZN(_16619_));
 AND2_X1 _36556_ (.A1(_11887_),
    .A2(_11886_),
    .ZN(_16598_));
 AND2_X1 _36557_ (.A1(_11888_),
    .A2(_11882_),
    .ZN(_16597_));
 AND2_X1 _36558_ (.A1(_11866_),
    .A2(_11879_),
    .ZN(_16605_));
 BUF_X2 _36559_ (.A(_11650_),
    .Z(_11889_));
 AND2_X1 _36560_ (.A1(_11889_),
    .A2(_11881_),
    .ZN(_16606_));
 AND2_X1 _36561_ (.A1(_11885_),
    .A2(_11880_),
    .ZN(_16607_));
 AND2_X1 _36562_ (.A1(_11853_),
    .A2(_11880_),
    .ZN(_17931_));
 AND2_X1 _36563_ (.A1(_11866_),
    .A2(_11886_),
    .ZN(_17930_));
 AND2_X1 _36564_ (.A1(_11865_),
    .A2(_11881_),
    .ZN(_17932_));
 AND2_X1 _36565_ (.A1(_11887_),
    .A2(_11686_),
    .ZN(_20880_));
 AND2_X1 _36566_ (.A1(_11860_),
    .A2(_11879_),
    .ZN(_17939_));
 NOR2_X1 _36567_ (.A1(_15313_),
    .A2(_18712_),
    .ZN(_17940_));
 BUF_X2 _36568_ (.A(_11662_),
    .Z(_11890_));
 AND2_X1 _36569_ (.A1(_11890_),
    .A2(_11882_),
    .ZN(_20882_));
 AND2_X1 _36570_ (.A1(_11865_),
    .A2(_11883_),
    .ZN(_20883_));
 AND2_X1 _36571_ (.A1(_11889_),
    .A2(_11685_),
    .ZN(_16677_));
 AND2_X1 _36572_ (.A1(_11866_),
    .A2(_11884_),
    .ZN(_16676_));
 AND2_X1 _36573_ (.A1(_11885_),
    .A2(_11686_),
    .ZN(_16675_));
 AND2_X1 _36574_ (.A1(_11885_),
    .A2(_11884_),
    .ZN(_16639_));
 AND2_X1 _36575_ (.A1(_11887_),
    .A2(_11685_),
    .ZN(_16640_));
 AND2_X1 _36576_ (.A1(_11889_),
    .A2(_11686_),
    .ZN(_16641_));
 AND2_X1 _36577_ (.A1(_11860_),
    .A2(_11881_),
    .ZN(_20877_));
 BUF_X2 _36578_ (.A(_11665_),
    .Z(_11891_));
 AND2_X1 _36579_ (.A1(_11891_),
    .A2(_11880_),
    .ZN(_20876_));
 AND2_X1 _36580_ (.A1(_11890_),
    .A2(_11886_),
    .ZN(_16643_));
 BUF_X1 _36581_ (.A(_11647_),
    .Z(_11892_));
 AND2_X1 _36582_ (.A1(_11892_),
    .A2(_11883_),
    .ZN(_16644_));
 AND2_X1 _36583_ (.A1(_11865_),
    .A2(_11882_),
    .ZN(_16645_));
 AND2_X1 _36584_ (.A1(_11892_),
    .A2(_11882_),
    .ZN(_16659_));
 AND2_X1 _36585_ (.A1(_11889_),
    .A2(_11884_),
    .ZN(_16658_));
 AND2_X1 _36586_ (.A1(_11885_),
    .A2(_11883_),
    .ZN(_16657_));
 AND2_X1 _36587_ (.A1(_11865_),
    .A2(_11886_),
    .ZN(_16662_));
 AND2_X1 _36588_ (.A1(_11860_),
    .A2(_11880_),
    .ZN(_16663_));
 AND2_X1 _36589_ (.A1(_11890_),
    .A2(_11881_),
    .ZN(_16664_));
 AND2_X1 _36590_ (.A1(_11857_),
    .A2(_11880_),
    .ZN(_18224_));
 BUF_X1 _36591_ (.A(_11656_),
    .Z(_11893_));
 AND2_X1 _36592_ (.A1(_11893_),
    .A2(_11886_),
    .ZN(_18223_));
 AND2_X1 _36593_ (.A1(_11891_),
    .A2(_11881_),
    .ZN(_18222_));
 AND2_X1 _36594_ (.A1(_11892_),
    .A2(_11686_),
    .ZN(_21054_));
 AND2_X1 _36595_ (.A1(_11885_),
    .A2(_11685_),
    .ZN(_21055_));
 AND2_X1 _36596_ (.A1(_11892_),
    .A2(_11685_),
    .ZN(_16680_));
 AND2_X1 _36597_ (.A1(_11890_),
    .A2(_11884_),
    .ZN(_16681_));
 BUF_X2 _36598_ (.A(_11659_),
    .Z(_11894_));
 AND2_X1 _36599_ (.A1(_11894_),
    .A2(_11686_),
    .ZN(_16682_));
 AND2_X1 _36600_ (.A1(_11890_),
    .A2(_11686_),
    .ZN(_21082_));
 AND2_X1 _36601_ (.A1(_11894_),
    .A2(_11685_),
    .ZN(_21081_));
 AND2_X1 _36602_ (.A1(_11893_),
    .A2(_11883_),
    .ZN(_20886_));
 AND2_X1 _36603_ (.A1(_11891_),
    .A2(_11882_),
    .ZN(_20885_));
 AND2_X1 _36604_ (.A1(_11857_),
    .A2(_11882_),
    .ZN(_18585_));
 AND2_X1 _36605_ (.A1(_11893_),
    .A2(_11884_),
    .ZN(_18586_));
 AND2_X1 _36606_ (.A1(_11891_),
    .A2(_11883_),
    .ZN(_18587_));
 BUF_X2 _36607_ (.A(a[89]),
    .Z(_11895_));
 AND2_X1 _36608_ (.A1(_11874_),
    .A2(_11895_),
    .ZN(_16737_));
 BUF_X2 _36609_ (.A(net220),
    .Z(_11896_));
 AND2_X1 _36610_ (.A1(_11837_),
    .A2(_11896_),
    .ZN(_16738_));
 BUF_X2 _36611_ (.A(net219),
    .Z(_11897_));
 AND2_X1 _36612_ (.A1(_11874_),
    .A2(_11897_),
    .ZN(_16749_));
 BUF_X2 _36613_ (.A(_11824_),
    .Z(_11898_));
 BUF_X2 _36614_ (.A(net218),
    .Z(_11899_));
 AND2_X1 _36615_ (.A1(_11898_),
    .A2(_11899_),
    .ZN(_16750_));
 AND2_X1 _36616_ (.A1(_11898_),
    .A2(_11897_),
    .ZN(_16747_));
 AND2_X1 _36617_ (.A1(_11841_),
    .A2(_11896_),
    .ZN(_18133_));
 INV_X2 _36618_ (.A(_11895_),
    .ZN(_18945_));
 NOR2_X1 _36619_ (.A1(_15964_),
    .A2(_18945_),
    .ZN(_18132_));
 AND2_X1 _36620_ (.A1(_11874_),
    .A2(_11899_),
    .ZN(_18141_));
 BUF_X2 _36621_ (.A(net217),
    .Z(_11900_));
 AND2_X1 _36622_ (.A1(_11898_),
    .A2(_11900_),
    .ZN(_18142_));
 AND2_X1 _36623_ (.A1(_11841_),
    .A2(_11897_),
    .ZN(_18136_));
 AND2_X1 _36624_ (.A1(_11845_),
    .A2(_11895_),
    .ZN(_18137_));
 AND2_X1 _36625_ (.A1(_11849_),
    .A2(_11896_),
    .ZN(_18138_));
 AND2_X1 _36626_ (.A1(_11848_),
    .A2(_11896_),
    .ZN(_16809_));
 AND2_X1 _36627_ (.A1(_11845_),
    .A2(_11899_),
    .ZN(_16808_));
 AND2_X1 _36628_ (.A1(_11842_),
    .A2(_11897_),
    .ZN(_16807_));
 BUF_X2 _36629_ (.A(net216),
    .Z(_11901_));
 AND2_X1 _36630_ (.A1(_11841_),
    .A2(_11901_),
    .ZN(_20891_));
 AND2_X1 _36631_ (.A1(_11849_),
    .A2(_11900_),
    .ZN(_20892_));
 BUF_X2 _36632_ (.A(net215),
    .Z(_11902_));
 AND2_X1 _36633_ (.A1(_11841_),
    .A2(_11902_),
    .ZN(_20893_));
 AND2_X1 _36634_ (.A1(_11849_),
    .A2(_11901_),
    .ZN(_20894_));
 AND2_X1 _36635_ (.A1(_11874_),
    .A2(_11902_),
    .ZN(_16754_));
 BUF_X2 _36636_ (.A(net214),
    .Z(_11903_));
 AND2_X1 _36637_ (.A1(_11898_),
    .A2(_11903_),
    .ZN(_16753_));
 AND2_X1 _36638_ (.A1(_11874_),
    .A2(_11903_),
    .ZN(_16803_));
 AND2_X1 _36639_ (.A1(_11898_),
    .A2(_11846_),
    .ZN(_16804_));
 AND2_X1 _36640_ (.A1(_11845_),
    .A2(_11897_),
    .ZN(_16769_));
 AND2_X1 _36641_ (.A1(_11841_),
    .A2(_11900_),
    .ZN(_16770_));
 AND2_X1 _36642_ (.A1(_11849_),
    .A2(_11899_),
    .ZN(_16771_));
 AND2_X1 _36643_ (.A1(_11874_),
    .A2(_11901_),
    .ZN(_16757_));
 AND2_X1 _36644_ (.A1(_11898_),
    .A2(_11902_),
    .ZN(_16758_));
 AND2_X1 _36645_ (.A1(_11842_),
    .A2(_11896_),
    .ZN(_16775_));
 NOR2_X1 _36646_ (.A1(_15915_),
    .A2(_18945_),
    .ZN(_16774_));
 AND2_X1 _36647_ (.A1(_11874_),
    .A2(_11900_),
    .ZN(_16782_));
 AND2_X1 _36648_ (.A1(_11898_),
    .A2(_11901_),
    .ZN(_16783_));
 AND2_X1 _36649_ (.A1(_11845_),
    .A2(_11896_),
    .ZN(_16790_));
 AND2_X1 _36650_ (.A1(_11841_),
    .A2(_11899_),
    .ZN(_16791_));
 AND2_X1 _36651_ (.A1(_11849_),
    .A2(_11897_),
    .ZN(_16792_));
 AND2_X1 _36652_ (.A1(_11898_),
    .A2(_11847_),
    .ZN(_20996_));
 AND2_X1 _36653_ (.A1(_11874_),
    .A2(_11846_),
    .ZN(_20995_));
 AND2_X1 _36654_ (.A1(_11848_),
    .A2(_11897_),
    .ZN(_17517_));
 AND2_X1 _36655_ (.A1(_11845_),
    .A2(_11900_),
    .ZN(_17518_));
 BUF_X1 _36656_ (.A(_11801_),
    .Z(_11904_));
 AND2_X1 _36657_ (.A1(_11904_),
    .A2(_11899_),
    .ZN(_17519_));
 AND2_X1 _36658_ (.A1(_11850_),
    .A2(_11896_),
    .ZN(_17523_));
 NOR2_X1 _36659_ (.A1(_15870_),
    .A2(_18945_),
    .ZN(_17522_));
 AND2_X1 _36660_ (.A1(_11851_),
    .A2(_11897_),
    .ZN(_16848_));
 AND2_X1 _36661_ (.A1(_11850_),
    .A2(_11900_),
    .ZN(_16849_));
 AND2_X1 _36662_ (.A1(_11852_),
    .A2(_11899_),
    .ZN(_16850_));
 AND2_X1 _36663_ (.A1(_11904_),
    .A2(_11902_),
    .ZN(_20898_));
 AND2_X1 _36664_ (.A1(_11848_),
    .A2(_11901_),
    .ZN(_20899_));
 AND2_X1 _36665_ (.A1(_11845_),
    .A2(_11903_),
    .ZN(_16825_));
 BUF_X2 _36666_ (.A(_11819_),
    .Z(_11905_));
 AND2_X1 _36667_ (.A1(_11905_),
    .A2(_11847_),
    .ZN(_16824_));
 AND2_X1 _36668_ (.A1(_11849_),
    .A2(_11846_),
    .ZN(_16826_));
 AND2_X1 _36669_ (.A1(_11849_),
    .A2(_11847_),
    .ZN(_20905_));
 CLKBUF_X3 _36670_ (.A(_11808_),
    .Z(_11906_));
 AND2_X1 _36671_ (.A1(_11906_),
    .A2(_11846_),
    .ZN(_20906_));
 AND2_X1 _36672_ (.A1(_11874_),
    .A2(_11847_),
    .ZN(_16833_));
 AND2_X1 _36673_ (.A1(_11849_),
    .A2(_11903_),
    .ZN(_16834_));
 AND2_X1 _36674_ (.A1(_11905_),
    .A2(_11846_),
    .ZN(_16835_));
 AND2_X1 _36675_ (.A1(_11850_),
    .A2(_11899_),
    .ZN(_20902_));
 AND2_X1 _36676_ (.A1(_11852_),
    .A2(_11897_),
    .ZN(_20903_));
 AND2_X1 _36677_ (.A1(_11848_),
    .A2(_11900_),
    .ZN(_16838_));
 AND2_X1 _36678_ (.A1(_11906_),
    .A2(_11902_),
    .ZN(_16839_));
 AND2_X1 _36679_ (.A1(_11904_),
    .A2(_11901_),
    .ZN(_16840_));
 AND2_X1 _36680_ (.A1(_11850_),
    .A2(_11901_),
    .ZN(_18428_));
 AND2_X1 _36681_ (.A1(_11904_),
    .A2(_11903_),
    .ZN(_18429_));
 AND2_X1 _36682_ (.A1(_11848_),
    .A2(_11902_),
    .ZN(_18430_));
 AND2_X1 _36683_ (.A1(_11850_),
    .A2(_11846_),
    .ZN(_20908_));
 BUF_X2 _36684_ (.A(_11800_),
    .Z(_11907_));
 AND2_X1 _36685_ (.A1(_11907_),
    .A2(_11847_),
    .ZN(_20909_));
 AND2_X1 _36686_ (.A1(_11852_),
    .A2(_11903_),
    .ZN(_18950_));
 AND2_X1 _36687_ (.A1(_11851_),
    .A2(_11902_),
    .ZN(_18949_));
 BUF_X2 _36688_ (.A(a[73]),
    .Z(_11908_));
 INV_X2 _36689_ (.A(_11908_),
    .ZN(_18898_));
 NOR2_X1 _36690_ (.A1(_18713_),
    .A2(_18898_),
    .ZN(_18420_));
 BUF_X2 _36691_ (.A(net204),
    .Z(_11909_));
 AND2_X1 _36692_ (.A1(_11889_),
    .A2(_11909_),
    .ZN(_16853_));
 NOR2_X1 _36693_ (.A1(_15196_),
    .A2(_18898_),
    .ZN(_16854_));
 BUF_X2 _36694_ (.A(net202),
    .Z(_11910_));
 AND2_X1 _36695_ (.A1(_11889_),
    .A2(_11910_),
    .ZN(_16897_));
 AND2_X1 _36696_ (.A1(_11892_),
    .A2(_11909_),
    .ZN(_16896_));
 BUF_X2 _36697_ (.A(net203),
    .Z(_11911_));
 AND2_X1 _36698_ (.A1(_11885_),
    .A2(_11911_),
    .ZN(_16895_));
 BUF_X2 _36699_ (.A(net200),
    .Z(_11912_));
 AND2_X1 _36700_ (.A1(_11887_),
    .A2(_11912_),
    .ZN(_16892_));
 BUF_X2 _36701_ (.A(net199),
    .Z(_11913_));
 AND2_X1 _36702_ (.A1(_11888_),
    .A2(_11913_),
    .ZN(_16893_));
 AND2_X1 _36703_ (.A1(_11887_),
    .A2(_11913_),
    .ZN(_16884_));
 BUF_X2 _36704_ (.A(net198),
    .Z(_11914_));
 AND2_X1 _36705_ (.A1(_11888_),
    .A2(_11914_),
    .ZN(_16885_));
 AND2_X1 _36706_ (.A1(_11892_),
    .A2(_11908_),
    .ZN(_16859_));
 AND2_X1 _36707_ (.A1(_11889_),
    .A2(_11911_),
    .ZN(_16858_));
 AND2_X1 _36708_ (.A1(_11885_),
    .A2(_11909_),
    .ZN(_16857_));
 AND2_X1 _36709_ (.A1(_11887_),
    .A2(_11910_),
    .ZN(_16862_));
 AND2_X1 _36710_ (.A1(_11888_),
    .A2(_11912_),
    .ZN(_16863_));
 AND2_X1 _36711_ (.A1(_11887_),
    .A2(_11911_),
    .ZN(_16872_));
 AND2_X1 _36712_ (.A1(_11888_),
    .A2(_11910_),
    .ZN(_16871_));
 AND2_X1 _36713_ (.A1(_11887_),
    .A2(_11914_),
    .ZN(_18078_));
 BUF_X2 _36714_ (.A(net197),
    .Z(_11915_));
 AND2_X1 _36715_ (.A1(_11888_),
    .A2(_11915_),
    .ZN(_18077_));
 AND2_X1 _36716_ (.A1(_11889_),
    .A2(_11913_),
    .ZN(_21044_));
 AND2_X1 _36717_ (.A1(_11885_),
    .A2(_11912_),
    .ZN(_21045_));
 AND2_X1 _36718_ (.A1(_11889_),
    .A2(_11912_),
    .ZN(_18088_));
 AND2_X1 _36719_ (.A1(_11892_),
    .A2(_11911_),
    .ZN(_18087_));
 AND2_X1 _36720_ (.A1(_11654_),
    .A2(_11910_),
    .ZN(_18086_));
 AND2_X1 _36721_ (.A1(_11894_),
    .A2(_11909_),
    .ZN(_18094_));
 NOR2_X1 _36722_ (.A1(_15238_),
    .A2(_18898_),
    .ZN(_18095_));
 AND2_X1 _36723_ (.A1(_11892_),
    .A2(_11913_),
    .ZN(_16910_));
 AND2_X1 _36724_ (.A1(_11889_),
    .A2(_11915_),
    .ZN(_16909_));
 AND2_X1 _36725_ (.A1(_11654_),
    .A2(_11914_),
    .ZN(_16908_));
 AND2_X1 _36726_ (.A1(_11888_),
    .A2(_11814_),
    .ZN(_20911_));
 AND2_X1 _36727_ (.A1(_11887_),
    .A2(_11813_),
    .ZN(_20912_));
 AND2_X1 _36728_ (.A1(_11893_),
    .A2(_11911_),
    .ZN(_16914_));
 AND2_X1 _36729_ (.A1(_11894_),
    .A2(_11912_),
    .ZN(_16913_));
 AND2_X1 _36730_ (.A1(_11890_),
    .A2(_11910_),
    .ZN(_16915_));
 AND2_X1 _36731_ (.A1(_11891_),
    .A2(_11911_),
    .ZN(_20918_));
 AND2_X1 _36732_ (.A1(_11893_),
    .A2(_11910_),
    .ZN(_20919_));
 AND2_X1 _36733_ (.A1(_11654_),
    .A2(_11915_),
    .ZN(_16951_));
 AND2_X1 _36734_ (.A1(_11645_),
    .A2(_11814_),
    .ZN(_16950_));
 AND2_X1 _36735_ (.A1(_11651_),
    .A2(_11813_),
    .ZN(_16949_));
 AND2_X1 _36736_ (.A1(_11892_),
    .A2(_11914_),
    .ZN(_16953_));
 AND2_X1 _36737_ (.A1(_11890_),
    .A2(_11912_),
    .ZN(_16954_));
 AND2_X1 _36738_ (.A1(_11894_),
    .A2(_11913_),
    .ZN(_16955_));
 AND2_X1 _36739_ (.A1(_11890_),
    .A2(_11911_),
    .ZN(_16922_));
 AND2_X1 _36740_ (.A1(_11892_),
    .A2(_11912_),
    .ZN(_16923_));
 AND2_X1 _36741_ (.A1(_11894_),
    .A2(_11910_),
    .ZN(_16924_));
 AND2_X1 _36742_ (.A1(_11651_),
    .A2(_11914_),
    .ZN(_20915_));
 AND2_X1 _36743_ (.A1(_11654_),
    .A2(_11913_),
    .ZN(_20914_));
 AND2_X1 _36744_ (.A1(_11645_),
    .A2(_11915_),
    .ZN(_16927_));
 AND2_X1 _36745_ (.A1(_11888_),
    .A2(_11813_),
    .ZN(_16928_));
 AND2_X1 _36746_ (.A1(_11893_),
    .A2(_11909_),
    .ZN(_16936_));
 NOR2_X1 _36747_ (.A1(_15313_),
    .A2(_18898_),
    .ZN(_16935_));
 AND2_X1 _36748_ (.A1(_11894_),
    .A2(_11914_),
    .ZN(_20998_));
 AND2_X1 _36749_ (.A1(_11890_),
    .A2(_11913_),
    .ZN(_20999_));
 AND2_X1 _36750_ (.A1(_11651_),
    .A2(_11814_),
    .ZN(_17558_));
 AND2_X1 _36751_ (.A1(_11648_),
    .A2(_11915_),
    .ZN(_17559_));
 AND2_X1 _36752_ (.A1(_11654_),
    .A2(_11813_),
    .ZN(_17557_));
 AND2_X1 _36753_ (.A1(_11648_),
    .A2(_11814_),
    .ZN(_16971_));
 AND2_X1 _36754_ (.A1(_11890_),
    .A2(_11915_),
    .ZN(_16973_));
 AND2_X1 _36755_ (.A1(_11894_),
    .A2(_11813_),
    .ZN(_16972_));
 AND2_X1 _36756_ (.A1(_11893_),
    .A2(_11913_),
    .ZN(_16958_));
 AND2_X1 _36757_ (.A1(_11894_),
    .A2(_11915_),
    .ZN(_16957_));
 AND2_X1 _36758_ (.A1(_11663_),
    .A2(_11914_),
    .ZN(_16959_));
 AND2_X1 _36759_ (.A1(_11891_),
    .A2(_11913_),
    .ZN(_21072_));
 AND2_X1 _36760_ (.A1(_11893_),
    .A2(_11914_),
    .ZN(_21073_));
 AND2_X1 _36761_ (.A1(_11654_),
    .A2(_11814_),
    .ZN(_20922_));
 AND2_X1 _36762_ (.A1(_11648_),
    .A2(_11813_),
    .ZN(_20921_));
 AND2_X1 _36763_ (.A1(_11894_),
    .A2(_11814_),
    .ZN(_21041_));
 AND2_X1 _36764_ (.A1(_11663_),
    .A2(_11813_),
    .ZN(_21042_));
 BUF_X1 _36765_ (.A(_11670_),
    .Z(_11916_));
 BUF_X2 _36766_ (.A(a[55]),
    .Z(_11917_));
 AND2_X1 _36767_ (.A1(_11916_),
    .A2(_11917_),
    .ZN(_16988_));
 BUF_X2 _36768_ (.A(net186),
    .Z(_11918_));
 AND2_X1 _36769_ (.A1(_11746_),
    .A2(_11918_),
    .ZN(_16989_));
 INV_X2 _36770_ (.A(_11917_),
    .ZN(_16975_));
 NOR2_X1 _36771_ (.A1(_18850_),
    .A2(_16975_),
    .ZN(_16985_));
 BUF_X2 _36772_ (.A(net187),
    .Z(_11919_));
 AND2_X1 _36773_ (.A1(_11768_),
    .A2(_11919_),
    .ZN(_18052_));
 BUF_X2 _36774_ (.A(a[57]),
    .Z(_11920_));
 INV_X2 _36775_ (.A(_11920_),
    .ZN(_18849_));
 NOR2_X1 _36776_ (.A1(_14944_),
    .A2(_18849_),
    .ZN(_18053_));
 AND2_X1 _36777_ (.A1(_11916_),
    .A2(_11918_),
    .ZN(_18061_));
 BUF_X2 _36778_ (.A(net185),
    .Z(_11921_));
 AND2_X1 _36779_ (.A1(_11746_),
    .A2(_11921_),
    .ZN(_18062_));
 AND2_X1 _36780_ (.A1(_11768_),
    .A2(_11917_),
    .ZN(_18058_));
 AND2_X1 _36781_ (.A1(_11756_),
    .A2(_11920_),
    .ZN(_18057_));
 AND2_X1 _36782_ (.A1(_11760_),
    .A2(_11919_),
    .ZN(_18056_));
 BUF_X2 _36783_ (.A(net184),
    .Z(_11922_));
 AND2_X1 _36784_ (.A1(_11768_),
    .A2(_11922_),
    .ZN(_20924_));
 AND2_X1 _36785_ (.A1(_11760_),
    .A2(_11921_),
    .ZN(_20925_));
 AND2_X1 _36786_ (.A1(_11760_),
    .A2(_11922_),
    .ZN(_20927_));
 BUF_X2 _36787_ (.A(net183),
    .Z(_11923_));
 AND2_X1 _36788_ (.A1(_11768_),
    .A2(_11923_),
    .ZN(_20926_));
 AND2_X1 _36789_ (.A1(_11916_),
    .A2(_11923_),
    .ZN(_16992_));
 BUF_X2 _36790_ (.A(net182),
    .Z(_11924_));
 AND2_X1 _36791_ (.A1(_11746_),
    .A2(_11924_),
    .ZN(_16993_));
 AND2_X1 _36792_ (.A1(_11756_),
    .A2(_11918_),
    .ZN(_17051_));
 BUF_X2 _36793_ (.A(_11692_),
    .Z(_11925_));
 AND2_X1 _36794_ (.A1(_11925_),
    .A2(_11919_),
    .ZN(_17052_));
 AND2_X1 _36795_ (.A1(_11759_),
    .A2(_11917_),
    .ZN(_17050_));
 AND2_X1 _36796_ (.A1(_11916_),
    .A2(_11924_),
    .ZN(_17038_));
 BUF_X2 _36797_ (.A(_11673_),
    .Z(_11926_));
 AND2_X1 _36798_ (.A1(_11926_),
    .A2(_11794_),
    .ZN(_17039_));
 AND2_X1 _36799_ (.A1(_11756_),
    .A2(_11917_),
    .ZN(_17008_));
 AND2_X1 _36800_ (.A1(_11768_),
    .A2(_11921_),
    .ZN(_17009_));
 AND2_X1 _36801_ (.A1(_11760_),
    .A2(_11918_),
    .ZN(_17010_));
 AND2_X1 _36802_ (.A1(_11916_),
    .A2(_11922_),
    .ZN(_16997_));
 AND2_X1 _36803_ (.A1(_11926_),
    .A2(_11923_),
    .ZN(_16996_));
 AND2_X1 _36804_ (.A1(_11759_),
    .A2(_11919_),
    .ZN(_17013_));
 NOR2_X1 _36805_ (.A1(_14888_),
    .A2(_18849_),
    .ZN(_17014_));
 AND2_X1 _36806_ (.A1(_11916_),
    .A2(_11921_),
    .ZN(_17022_));
 AND2_X1 _36807_ (.A1(_11926_),
    .A2(_11922_),
    .ZN(_17021_));
 AND2_X1 _36808_ (.A1(_11768_),
    .A2(_11918_),
    .ZN(_17029_));
 AND2_X1 _36809_ (.A1(_11756_),
    .A2(_11919_),
    .ZN(_17030_));
 NOR2_X1 _36810_ (.A1(_14944_),
    .A2(_16975_),
    .ZN(_17031_));
 AND2_X1 _36811_ (.A1(_11926_),
    .A2(_11795_),
    .ZN(_20929_));
 AND2_X1 _36812_ (.A1(_11916_),
    .A2(_11794_),
    .ZN(_20928_));
 NOR2_X1 _36813_ (.A1(_14888_),
    .A2(_16975_),
    .ZN(_17589_));
 AND2_X1 _36814_ (.A1(_11756_),
    .A2(_11921_),
    .ZN(_17590_));
 AND2_X1 _36815_ (.A1(_11759_),
    .A2(_11918_),
    .ZN(_17591_));
 AND2_X1 _36816_ (.A1(_11741_),
    .A2(_11919_),
    .ZN(_17594_));
 NOR2_X1 _36817_ (.A1(_14841_),
    .A2(_18849_),
    .ZN(_17595_));
 AND2_X1 _36818_ (.A1(_11756_),
    .A2(_11922_),
    .ZN(_17060_));
 AND2_X1 _36819_ (.A1(_11768_),
    .A2(_11924_),
    .ZN(_17059_));
 AND2_X1 _36820_ (.A1(_11760_),
    .A2(_11923_),
    .ZN(_17058_));
 AND2_X1 _36821_ (.A1(_11741_),
    .A2(_11917_),
    .ZN(_17068_));
 AND2_X1 _36822_ (.A1(_11759_),
    .A2(_11921_),
    .ZN(_17069_));
 AND2_X1 _36823_ (.A1(_11925_),
    .A2(_11918_),
    .ZN(_17070_));
 AND2_X1 _36824_ (.A1(_11760_),
    .A2(_11924_),
    .ZN(_17083_));
 AND2_X1 _36825_ (.A1(_11916_),
    .A2(_11795_),
    .ZN(_17082_));
 AND2_X1 _36826_ (.A1(_11768_),
    .A2(_11794_),
    .ZN(_17084_));
 NOR2_X1 _36827_ (.A1(_14841_),
    .A2(_16975_),
    .ZN(_20932_));
 BUF_X2 _36828_ (.A(_11690_),
    .Z(_11927_));
 AND2_X1 _36829_ (.A1(_11927_),
    .A2(_11918_),
    .ZN(_20933_));
 AND2_X1 _36830_ (.A1(_11925_),
    .A2(_11921_),
    .ZN(_17088_));
 BUF_X1 _36831_ (.A(_11683_),
    .Z(_11928_));
 AND2_X1 _36832_ (.A1(_11928_),
    .A2(_11923_),
    .ZN(_17087_));
 AND2_X1 _36833_ (.A1(_11759_),
    .A2(_11922_),
    .ZN(_17086_));
 AND2_X1 _36834_ (.A1(_11759_),
    .A2(_11923_),
    .ZN(_20935_));
 AND2_X1 _36835_ (.A1(_11925_),
    .A2(_11922_),
    .ZN(_20936_));
 AND2_X1 _36836_ (.A1(_11928_),
    .A2(_11924_),
    .ZN(_17101_));
 AND2_X1 _36837_ (.A1(_11768_),
    .A2(_11795_),
    .ZN(_17100_));
 BUF_X2 _36838_ (.A(_11680_),
    .Z(_11929_));
 AND2_X1 _36839_ (.A1(_11929_),
    .A2(_11794_),
    .ZN(_17099_));
 AND2_X1 _36840_ (.A1(_11927_),
    .A2(_11921_),
    .ZN(_18033_));
 AND2_X1 _36841_ (.A1(_11781_),
    .A2(_11917_),
    .ZN(_18032_));
 AND2_X1 _36842_ (.A1(_11732_),
    .A2(_11918_),
    .ZN(_18034_));
 AND2_X1 _36843_ (.A1(_11929_),
    .A2(_11795_),
    .ZN(_21039_));
 AND2_X1 _36844_ (.A1(_11928_),
    .A2(_11794_),
    .ZN(_21038_));
 AND2_X1 _36845_ (.A1(_11927_),
    .A2(_11923_),
    .ZN(_20937_));
 AND2_X1 _36846_ (.A1(_11732_),
    .A2(_11922_),
    .ZN(_20938_));
 AND2_X1 _36847_ (.A1(_11925_),
    .A2(_11924_),
    .ZN(_17106_));
 AND2_X1 _36848_ (.A1(_11928_),
    .A2(_11795_),
    .ZN(_17105_));
 BUF_X2 _36849_ (.A(_11725_),
    .Z(_11930_));
 AND2_X1 _36850_ (.A1(_11930_),
    .A2(_11794_),
    .ZN(_17104_));
 AND2_X1 _36851_ (.A1(_11930_),
    .A2(_11795_),
    .ZN(_21079_));
 AND2_X1 _36852_ (.A1(_11925_),
    .A2(_11794_),
    .ZN(_21080_));
 AND2_X1 _36853_ (.A1(_11927_),
    .A2(_11924_),
    .ZN(_18538_));
 AND2_X1 _36854_ (.A1(_11781_),
    .A2(_11922_),
    .ZN(_18537_));
 BUF_X1 _36855_ (.A(_11688_),
    .Z(_11931_));
 AND2_X1 _36856_ (.A1(_11931_),
    .A2(_11923_),
    .ZN(_18536_));
 BUF_X2 _36857_ (.A(net170),
    .Z(_11932_));
 AND2_X1 _36858_ (.A1(_11792_),
    .A2(_11932_),
    .ZN(_17125_));
 BUF_X2 _36859_ (.A(net169),
    .Z(_11933_));
 AND2_X1 _36860_ (.A1(_11793_),
    .A2(_11933_),
    .ZN(_17126_));
 AND2_X1 _36861_ (.A1(_11793_),
    .A2(_11932_),
    .ZN(_17123_));
 BUF_X2 _36862_ (.A(a[41]),
    .Z(_11934_));
 AND2_X1 _36863_ (.A1(_11792_),
    .A2(_11934_),
    .ZN(_17118_));
 BUF_X2 _36864_ (.A(net172),
    .Z(_11935_));
 AND2_X1 _36865_ (.A1(_11793_),
    .A2(_11935_),
    .ZN(_17119_));
 AND2_X1 _36866_ (.A1(_11790_),
    .A2(_11935_),
    .ZN(_17605_));
 INV_X2 _36867_ (.A(_11934_),
    .ZN(_18804_));
 NOR2_X1 _36868_ (.A1(_15651_),
    .A2(_18804_),
    .ZN(_17606_));
 AND2_X1 _36869_ (.A1(_11792_),
    .A2(_11933_),
    .ZN(_17615_));
 BUF_X2 _36870_ (.A(net168),
    .Z(_11936_));
 AND2_X1 _36871_ (.A1(_11793_),
    .A2(_11936_),
    .ZN(_17614_));
 AND2_X1 _36872_ (.A1(_11791_),
    .A2(_11934_),
    .ZN(_17609_));
 AND2_X1 _36873_ (.A1(_11790_),
    .A2(_11932_),
    .ZN(_17610_));
 AND2_X1 _36874_ (.A1(_11796_),
    .A2(_11935_),
    .ZN(_17611_));
 BUF_X2 _36875_ (.A(net167),
    .Z(_11937_));
 AND2_X1 _36876_ (.A1(_11792_),
    .A2(_11937_),
    .ZN(_17146_));
 BUF_X2 _36877_ (.A(net166),
    .Z(_11938_));
 AND2_X1 _36878_ (.A1(_11793_),
    .A2(_11938_),
    .ZN(_17147_));
 AND2_X1 _36879_ (.A1(_11792_),
    .A2(_11936_),
    .ZN(_17134_));
 AND2_X1 _36880_ (.A1(_11793_),
    .A2(_11937_),
    .ZN(_17133_));
 AND2_X1 _36881_ (.A1(_11790_),
    .A2(_11933_),
    .ZN(_17138_));
 AND2_X1 _36882_ (.A1(_11791_),
    .A2(_11935_),
    .ZN(_17137_));
 AND2_X1 _36883_ (.A1(_11796_),
    .A2(_11932_),
    .ZN(_17139_));
 AND2_X1 _36884_ (.A1(_11792_),
    .A2(_11938_),
    .ZN(_17155_));
 BUF_X2 _36885_ (.A(_11712_),
    .Z(_11939_));
 BUF_X2 _36886_ (.A(net165),
    .Z(_11940_));
 AND2_X1 _36887_ (.A1(_11939_),
    .A2(_11940_),
    .ZN(_17156_));
 AND2_X1 _36888_ (.A1(_11796_),
    .A2(_11936_),
    .ZN(_20940_));
 AND2_X1 _36889_ (.A1(_11790_),
    .A2(_11937_),
    .ZN(_20941_));
 BUF_X2 _36890_ (.A(_11705_),
    .Z(_11941_));
 AND2_X1 _36891_ (.A1(_11941_),
    .A2(_11936_),
    .ZN(_17159_));
 AND2_X1 _36892_ (.A1(_11791_),
    .A2(_11932_),
    .ZN(_17160_));
 AND2_X1 _36893_ (.A1(_11796_),
    .A2(_11933_),
    .ZN(_17161_));
 AND2_X1 _36894_ (.A1(_11786_),
    .A2(_11935_),
    .ZN(_17167_));
 NOR2_X1 _36895_ (.A1(_15412_),
    .A2(_18804_),
    .ZN(_17168_));
 AND2_X1 _36896_ (.A1(_11791_),
    .A2(_11933_),
    .ZN(_17185_));
 AND2_X1 _36897_ (.A1(_11787_),
    .A2(_11935_),
    .ZN(_17184_));
 BUF_X2 _36898_ (.A(_11700_),
    .Z(_11942_));
 AND2_X1 _36899_ (.A1(_11942_),
    .A2(_11932_),
    .ZN(_17183_));
 AND2_X1 _36900_ (.A1(_11796_),
    .A2(_11937_),
    .ZN(_20944_));
 AND2_X1 _36901_ (.A1(_11941_),
    .A2(_11938_),
    .ZN(_20945_));
 BUF_X1 _36902_ (.A(_11703_),
    .Z(_11943_));
 AND2_X1 _36903_ (.A1(_11943_),
    .A2(_11940_),
    .ZN(_17175_));
 AND2_X1 _36904_ (.A1(_11939_),
    .A2(_11773_),
    .ZN(_17176_));
 AND2_X1 _36905_ (.A1(_11787_),
    .A2(_11932_),
    .ZN(_18010_));
 BUF_X1 _36906_ (.A(_11697_),
    .Z(_11944_));
 AND2_X1 _36907_ (.A1(_11944_),
    .A2(_11936_),
    .ZN(_18009_));
 AND2_X1 _36908_ (.A1(_11942_),
    .A2(_11933_),
    .ZN(_18008_));
 AND2_X1 _36909_ (.A1(_11939_),
    .A2(_11771_),
    .ZN(_20946_));
 AND2_X1 _36910_ (.A1(_11943_),
    .A2(_11773_),
    .ZN(_20947_));
 AND2_X1 _36911_ (.A1(_11782_),
    .A2(_11935_),
    .ZN(_18018_));
 NOR2_X1 _36912_ (.A1(_14677_),
    .A2(_18804_),
    .ZN(_18017_));
 AND2_X1 _36913_ (.A1(_11944_),
    .A2(_11937_),
    .ZN(_17195_));
 AND2_X1 _36914_ (.A1(_11941_),
    .A2(_11940_),
    .ZN(_17196_));
 AND2_X1 _36915_ (.A1(_11796_),
    .A2(_11938_),
    .ZN(_17197_));
 AND2_X1 _36916_ (.A1(_11942_),
    .A2(_11936_),
    .ZN(_17205_));
 AND2_X1 _36917_ (.A1(_11782_),
    .A2(_11932_),
    .ZN(_17206_));
 AND2_X1 _36918_ (.A1(_11787_),
    .A2(_11933_),
    .ZN(_17207_));
 AND2_X1 _36919_ (.A1(_11782_),
    .A2(_11933_),
    .ZN(_20952_));
 AND2_X1 _36920_ (.A1(_11772_),
    .A2(_11932_),
    .ZN(_20951_));
 AND2_X1 _36921_ (.A1(_11796_),
    .A2(_11940_),
    .ZN(_17221_));
 AND2_X1 _36922_ (.A1(_11943_),
    .A2(_11771_),
    .ZN(_17220_));
 AND2_X1 _36923_ (.A1(_11941_),
    .A2(_11773_),
    .ZN(_17219_));
 BUF_X2 _36924_ (.A(_11695_),
    .Z(_11945_));
 AND2_X1 _36925_ (.A1(_11945_),
    .A2(_11936_),
    .ZN(_17224_));
 AND2_X1 _36926_ (.A1(_11944_),
    .A2(_11938_),
    .ZN(_17225_));
 AND2_X1 _36927_ (.A1(_11942_),
    .A2(_11937_),
    .ZN(_17226_));
 AND2_X1 _36928_ (.A1(_11942_),
    .A2(_11938_),
    .ZN(_20955_));
 AND2_X1 _36929_ (.A1(_11945_),
    .A2(_11937_),
    .ZN(_20954_));
 AND2_X1 _36930_ (.A1(_11944_),
    .A2(_11940_),
    .ZN(_17237_));
 AND2_X1 _36931_ (.A1(_11941_),
    .A2(_11771_),
    .ZN(_17238_));
 AND2_X1 _36932_ (.A1(_11796_),
    .A2(_11773_),
    .ZN(_17239_));
 BUF_X1 _36933_ (.A(_11776_),
    .Z(_11946_));
 AND2_X1 _36934_ (.A1(_11946_),
    .A2(_11932_),
    .ZN(_17987_));
 AND2_X1 _36935_ (.A1(_11782_),
    .A2(_11936_),
    .ZN(_17986_));
 AND2_X1 _36936_ (.A1(_11772_),
    .A2(_11933_),
    .ZN(_17985_));
 AND2_X1 _36937_ (.A1(_11796_),
    .A2(_11771_),
    .ZN(_21034_));
 AND2_X1 _36938_ (.A1(_11944_),
    .A2(_11773_),
    .ZN(_21035_));
 AND2_X1 _36939_ (.A1(_11772_),
    .A2(_11937_),
    .ZN(_20956_));
 AND2_X1 _36940_ (.A1(_11782_),
    .A2(_11938_),
    .ZN(_20957_));
 AND2_X1 _36941_ (.A1(_11944_),
    .A2(_11771_),
    .ZN(_17242_));
 AND2_X1 _36942_ (.A1(_11945_),
    .A2(_11940_),
    .ZN(_17244_));
 AND2_X1 _36943_ (.A1(_11942_),
    .A2(_11773_),
    .ZN(_17243_));
 AND2_X1 _36944_ (.A1(_11942_),
    .A2(_11771_),
    .ZN(_21077_));
 AND2_X1 _36945_ (.A1(_11945_),
    .A2(_11773_),
    .ZN(_21078_));
 BUF_X1 _36946_ (.A(_11715_),
    .Z(_11947_));
 AND2_X1 _36947_ (.A1(_11947_),
    .A2(_11940_),
    .ZN(_18487_));
 AND2_X1 _36948_ (.A1(_11946_),
    .A2(_11937_),
    .ZN(_18488_));
 AND2_X1 _36949_ (.A1(_11873_),
    .A2(_11938_),
    .ZN(_18489_));
 BUF_X2 _36950_ (.A(net89),
    .Z(_11948_));
 AND2_X1 _36951_ (.A1(_11812_),
    .A2(_11948_),
    .ZN(_17258_));
 AND2_X1 _36952_ (.A1(_11764_),
    .A2(_11821_),
    .ZN(_17257_));
 AND2_X1 _36953_ (.A1(_11767_),
    .A2(_11820_),
    .ZN(_17259_));
 BUF_X2 _36954_ (.A(a[23]),
    .Z(_11949_));
 INV_X2 _36955_ (.A(_11949_),
    .ZN(_17348_));
 NOR2_X1 _36956_ (.A1(_15870_),
    .A2(_17348_),
    .ZN(_20960_));
 BUF_X2 _36957_ (.A(net131),
    .Z(_11950_));
 AND2_X1 _36958_ (.A1(_11850_),
    .A2(_11950_),
    .ZN(_20961_));
 BUF_X2 _36959_ (.A(net99),
    .Z(_11951_));
 AND2_X1 _36960_ (.A1(_11906_),
    .A2(_11951_),
    .ZN(_17263_));
 BUF_X2 _36961_ (.A(net120),
    .Z(_11952_));
 AND2_X1 _36962_ (.A1(_11907_),
    .A2(_11952_),
    .ZN(_17262_));
 BUF_X2 _36963_ (.A(net110),
    .Z(_11953_));
 AND2_X1 _36964_ (.A1(_11904_),
    .A2(_11953_),
    .ZN(_17261_));
 AND2_X1 _36965_ (.A1(_11904_),
    .A2(_11951_),
    .ZN(_20967_));
 AND2_X1 _36966_ (.A1(_11907_),
    .A2(_11953_),
    .ZN(_20968_));
 AND2_X1 _36967_ (.A1(_11906_),
    .A2(_11948_),
    .ZN(_17295_));
 AND2_X1 _36968_ (.A1(_11764_),
    .A2(_11820_),
    .ZN(_17294_));
 AND2_X1 _36969_ (.A1(_11767_),
    .A2(_11811_),
    .ZN(_17293_));
 AND2_X1 _36970_ (.A1(_11905_),
    .A2(_11948_),
    .ZN(_17270_));
 AND2_X1 _36971_ (.A1(_11906_),
    .A2(_11953_),
    .ZN(_17271_));
 AND2_X1 _36972_ (.A1(_11812_),
    .A2(_11951_),
    .ZN(_17272_));
 AND2_X1 _36973_ (.A1(_11764_),
    .A2(_11824_),
    .ZN(_20963_));
 AND2_X1 _36974_ (.A1(_11767_),
    .A2(_11821_),
    .ZN(_20964_));
 AND2_X1 _36975_ (.A1(_11904_),
    .A2(_11952_),
    .ZN(_17281_));
 BUF_X1 _36976_ (.A(_11762_),
    .Z(_11954_));
 AND2_X1 _36977_ (.A1(_11954_),
    .A2(_11949_),
    .ZN(_17280_));
 AND2_X1 _36978_ (.A1(_11907_),
    .A2(_11950_),
    .ZN(_17282_));
 AND2_X1 _36979_ (.A1(_11954_),
    .A2(_11952_),
    .ZN(_17365_));
 AND2_X1 _36980_ (.A1(_11851_),
    .A2(_11949_),
    .ZN(_17366_));
 AND2_X1 _36981_ (.A1(_11852_),
    .A2(_11950_),
    .ZN(_17367_));
 AND2_X1 _36982_ (.A1(_11764_),
    .A2(_11811_),
    .ZN(_20976_));
 AND2_X1 _36983_ (.A1(_11767_),
    .A2(_11809_),
    .ZN(_20977_));
 AND2_X1 _36984_ (.A1(_11812_),
    .A2(_11953_),
    .ZN(_20970_));
 AND2_X1 _36985_ (.A1(_11905_),
    .A2(_11951_),
    .ZN(_20969_));
 AND2_X1 _36986_ (.A1(_11822_),
    .A2(_11948_),
    .ZN(_17298_));
 AND2_X1 _36987_ (.A1(_11767_),
    .A2(_11824_),
    .ZN(_17299_));
 NOR2_X1 _36988_ (.A1(_15915_),
    .A2(_17348_),
    .ZN(_17313_));
 AND2_X1 _36989_ (.A1(_11906_),
    .A2(_11952_),
    .ZN(_17312_));
 AND2_X1 _36990_ (.A1(_11904_),
    .A2(_11950_),
    .ZN(_17311_));
 BUF_X2 _36991_ (.A(net149),
    .Z(_11955_));
 AND2_X1 _36992_ (.A1(_11954_),
    .A2(_11955_),
    .ZN(_17316_));
 BUF_X2 _36993_ (.A(a[25]),
    .Z(_11956_));
 INV_X2 _36994_ (.A(_11956_),
    .ZN(_18756_));
 NOR2_X1 _36995_ (.A1(_15870_),
    .A2(_18756_),
    .ZN(_17317_));
 AND2_X1 _36996_ (.A1(_11905_),
    .A2(_11953_),
    .ZN(_20972_));
 AND2_X1 _36997_ (.A1(_11812_),
    .A2(_11952_),
    .ZN(_20973_));
 AND2_X1 _36998_ (.A1(_11822_),
    .A2(_11951_),
    .ZN(_17325_));
 AND2_X1 _36999_ (.A1(_11898_),
    .A2(_11948_),
    .ZN(_17324_));
 AND2_X1 _37000_ (.A1(_11907_),
    .A2(_11955_),
    .ZN(_17332_));
 AND2_X1 _37001_ (.A1(_11906_),
    .A2(_11950_),
    .ZN(_17333_));
 AND2_X1 _37002_ (.A1(_11904_),
    .A2(_11949_),
    .ZN(_17334_));
 AND2_X1 _37003_ (.A1(_11822_),
    .A2(_11949_),
    .ZN(_17361_));
 AND2_X1 _37004_ (.A1(_11898_),
    .A2(_11950_),
    .ZN(_17362_));
 NOR2_X1 _37005_ (.A1(_18757_),
    .A2(_17348_),
    .ZN(_17358_));
 AND2_X1 _37006_ (.A1(_11905_),
    .A2(_11955_),
    .ZN(_17389_));
 NOR2_X1 _37007_ (.A1(_15964_),
    .A2(_18756_),
    .ZN(_17390_));
 AND2_X1 _37008_ (.A1(_11822_),
    .A2(_11950_),
    .ZN(_17398_));
 AND2_X1 _37009_ (.A1(_11825_),
    .A2(_11952_),
    .ZN(_17399_));
 AND2_X1 _37010_ (.A1(_11906_),
    .A2(_11956_),
    .ZN(_17395_));
 AND2_X1 _37011_ (.A1(_11905_),
    .A2(_11949_),
    .ZN(_17394_));
 AND2_X1 _37012_ (.A1(_11812_),
    .A2(_11955_),
    .ZN(_17393_));
 AND2_X1 _37013_ (.A1(_11954_),
    .A2(_11767_),
    .ZN(_20974_));
 AND2_X1 _37014_ (.A1(_11764_),
    .A2(_11800_),
    .ZN(_20975_));
 AND2_X1 _37015_ (.A1(_11852_),
    .A2(_11948_),
    .ZN(_18762_));
 AND2_X1 _37016_ (.A1(_11851_),
    .A2(_11951_),
    .ZN(_18761_));
 AND2_X1 _37017_ (.A1(_11904_),
    .A2(_11948_),
    .ZN(_17380_));
 AND2_X1 _37018_ (.A1(_11954_),
    .A2(_11953_),
    .ZN(_17379_));
 AND2_X1 _37019_ (.A1(_11907_),
    .A2(_11951_),
    .ZN(_17381_));
 AND2_X1 _37020_ (.A1(_11764_),
    .A2(_11809_),
    .ZN(_17630_));
 AND2_X1 _37021_ (.A1(_11907_),
    .A2(_11948_),
    .ZN(_17631_));
 AND2_X1 _37022_ (.A1(_11767_),
    .A2(_11802_),
    .ZN(_17632_));
 AND2_X1 _37023_ (.A1(_11852_),
    .A2(_11953_),
    .ZN(_21002_));
 AND2_X1 _37024_ (.A1(_11954_),
    .A2(_11951_),
    .ZN(_21001_));
 AND2_X1 _37025_ (.A1(_11905_),
    .A2(_11950_),
    .ZN(_17422_));
 AND2_X1 _37026_ (.A1(_11906_),
    .A2(_11955_),
    .ZN(_17423_));
 NOR2_X1 _37027_ (.A1(_15964_),
    .A2(_17348_),
    .ZN(_17424_));
 AND2_X1 _37028_ (.A1(_11822_),
    .A2(_11952_),
    .ZN(_17415_));
 AND2_X1 _37029_ (.A1(_11825_),
    .A2(_11953_),
    .ZN(_17416_));
 AND2_X1 _37030_ (.A1(_11822_),
    .A2(_11953_),
    .ZN(_17412_));
 AND2_X1 _37031_ (.A1(_11825_),
    .A2(_11951_),
    .ZN(_17411_));
 AND2_X1 _37032_ (.A1(_11905_),
    .A2(_11952_),
    .ZN(_17961_));
 AND2_X1 _37033_ (.A1(_11906_),
    .A2(_11949_),
    .ZN(_17962_));
 AND2_X1 _37034_ (.A1(_11812_),
    .A2(_11950_),
    .ZN(_17963_));
 AND2_X1 _37035_ (.A1(_11802_),
    .A2(_11955_),
    .ZN(_17966_));
 NOR2_X1 _37036_ (.A1(_15915_),
    .A2(_18756_),
    .ZN(_17967_));
 BUF_X2 _37037_ (.A(net2),
    .Z(_11957_));
 AND2_X1 _37038_ (.A1(_11946_),
    .A2(_11957_),
    .ZN(_17428_));
 BUF_X2 _37039_ (.A(net230),
    .Z(_11958_));
 AND2_X1 _37040_ (.A1(_11947_),
    .A2(_11958_),
    .ZN(_17427_));
 BUF_X2 _37041_ (.A(net231),
    .Z(_11959_));
 AND2_X1 _37042_ (.A1(_11873_),
    .A2(_11959_),
    .ZN(_17426_));
 AND2_X1 _37043_ (.A1(_11942_),
    .A2(_11872_),
    .ZN(_20979_));
 AND2_X1 _37044_ (.A1(_11945_),
    .A2(_11871_),
    .ZN(_20980_));
 AND2_X1 _37045_ (.A1(_11945_),
    .A2(_11872_),
    .ZN(_21063_));
 AND2_X1 _37046_ (.A1(_11947_),
    .A2(_11871_),
    .ZN(_21064_));
 BUF_X2 _37047_ (.A(net15),
    .Z(_11960_));
 AND2_X1 _37048_ (.A1(_11925_),
    .A2(_11960_),
    .ZN(_17433_));
 AND2_X1 _37049_ (.A1(_11928_),
    .A2(_11876_),
    .ZN(_17432_));
 AND2_X1 _37050_ (.A1(_11930_),
    .A2(_11877_),
    .ZN(_17431_));
 AND2_X1 _37051_ (.A1(_11930_),
    .A2(_11876_),
    .ZN(_21068_));
 AND2_X1 _37052_ (.A1(_11925_),
    .A2(_11877_),
    .ZN(_21069_));
 BUF_X2 _37053_ (.A(net17),
    .Z(_11961_));
 AND2_X1 _37054_ (.A1(_11931_),
    .A2(_11961_),
    .ZN(_20983_));
 BUF_X2 _37055_ (.A(net16),
    .Z(_11962_));
 AND2_X1 _37056_ (.A1(_11927_),
    .A2(_11962_),
    .ZN(_20984_));
 AND2_X1 _37057_ (.A1(_11927_),
    .A2(_11960_),
    .ZN(_18324_));
 AND2_X1 _37058_ (.A1(_11781_),
    .A2(_11961_),
    .ZN(_18323_));
 AND2_X1 _37059_ (.A1(_11931_),
    .A2(_11962_),
    .ZN(_18322_));
 BUF_X2 _37060_ (.A(net5),
    .Z(_11963_));
 AND2_X1 _37061_ (.A1(_11945_),
    .A2(_11963_),
    .ZN(_17454_));
 BUF_X2 _37062_ (.A(net4),
    .Z(_11964_));
 AND2_X1 _37063_ (.A1(_11944_),
    .A2(_11964_),
    .ZN(_17455_));
 CLKBUF_X2 _37064_ (.A(a[103]),
    .Z(_11965_));
 AND2_X1 _37065_ (.A1(_11942_),
    .A2(_11965_),
    .ZN(_17456_));
 BUF_X2 _37066_ (.A(net3),
    .Z(_11966_));
 AND2_X1 _37067_ (.A1(_11709_),
    .A2(_11966_),
    .ZN(_20987_));
 AND2_X1 _37068_ (.A1(_11941_),
    .A2(_11957_),
    .ZN(_20986_));
 AND2_X1 _37069_ (.A1(_11941_),
    .A2(_11959_),
    .ZN(_20989_));
 AND2_X1 _37070_ (.A1(_11709_),
    .A2(_11957_),
    .ZN(_20988_));
 AND2_X1 _37071_ (.A1(_11943_),
    .A2(_11959_),
    .ZN(_17441_));
 AND2_X1 _37072_ (.A1(_11939_),
    .A2(_11958_),
    .ZN(_17442_));
 AND2_X1 _37073_ (.A1(_11943_),
    .A2(_11958_),
    .ZN(_17451_));
 AND2_X1 _37074_ (.A1(_11939_),
    .A2(_11871_),
    .ZN(_17450_));
 INV_X1 _37075_ (.A(_11965_),
    .ZN(_18314_));
 NOR2_X1 _37076_ (.A1(_15412_),
    .A2(_18314_),
    .ZN(_17497_));
 AND2_X1 _37077_ (.A1(_11944_),
    .A2(_11966_),
    .ZN(_17496_));
 AND2_X1 _37078_ (.A1(_11942_),
    .A2(_11964_),
    .ZN(_17495_));
 AND2_X1 _37079_ (.A1(_11939_),
    .A2(_11872_),
    .ZN(_20992_));
 AND2_X1 _37080_ (.A1(_11943_),
    .A2(_11871_),
    .ZN(_20993_));
 AND2_X1 _37081_ (.A1(_11947_),
    .A2(_11963_),
    .ZN(_17505_));
 BUF_X2 _37082_ (.A(a[105]),
    .Z(_11967_));
 INV_X2 _37083_ (.A(_11967_),
    .ZN(_18987_));
 NOR2_X1 _37084_ (.A1(_14677_),
    .A2(_18987_),
    .ZN(_17504_));
 AND2_X1 _37085_ (.A1(_11941_),
    .A2(_11966_),
    .ZN(_17471_));
 AND2_X1 _37086_ (.A1(_11944_),
    .A2(_11965_),
    .ZN(_17470_));
 AND2_X1 _37087_ (.A1(_11709_),
    .A2(_11964_),
    .ZN(_17472_));
 AND2_X1 _37088_ (.A1(_11943_),
    .A2(_11957_),
    .ZN(_17475_));
 AND2_X1 _37089_ (.A1(_11939_),
    .A2(_11959_),
    .ZN(_17476_));
 AND2_X1 _37090_ (.A1(_11701_),
    .A2(_11963_),
    .ZN(_17482_));
 NOR2_X1 _37091_ (.A1(_15412_),
    .A2(_18987_),
    .ZN(_17483_));
 AND2_X1 _37092_ (.A1(_11944_),
    .A2(_11957_),
    .ZN(_17872_));
 AND2_X1 _37093_ (.A1(_11941_),
    .A2(_11958_),
    .ZN(_17871_));
 AND2_X1 _37094_ (.A1(_11709_),
    .A2(_11959_),
    .ZN(_17870_));
 AND2_X1 _37095_ (.A1(_11701_),
    .A2(_11966_),
    .ZN(_17876_));
 AND2_X1 _37096_ (.A1(_11947_),
    .A2(_11965_),
    .ZN(_17875_));
 AND2_X1 _37097_ (.A1(_11945_),
    .A2(_11964_),
    .ZN(_17877_));
 AND2_X1 _37098_ (.A1(_11905_),
    .A2(_11903_),
    .ZN(_17539_));
 AND2_X1 _37099_ (.A1(_11809_),
    .A2(_11901_),
    .ZN(_17538_));
 AND2_X1 _37100_ (.A1(_11812_),
    .A2(_11902_),
    .ZN(_17540_));
 AND2_X1 _37101_ (.A1(_11802_),
    .A2(_11900_),
    .ZN(_17548_));
 AND2_X1 _37102_ (.A1(_11954_),
    .A2(_11897_),
    .ZN(_17549_));
 AND2_X1 _37103_ (.A1(_11907_),
    .A2(_11899_),
    .ZN(_17547_));
 AND2_X1 _37104_ (.A1(_11857_),
    .A2(_11911_),
    .ZN(_17573_));
 AND2_X1 _37105_ (.A1(_11893_),
    .A2(_11912_),
    .ZN(_17572_));
 AND2_X1 _37106_ (.A1(_11891_),
    .A2(_11910_),
    .ZN(_17571_));
 AND2_X1 _37107_ (.A1(_11764_),
    .A2(_11802_),
    .ZN(_21083_));
 AND2_X1 _37108_ (.A1(_11767_),
    .A2(_11800_),
    .ZN(_21084_));
 AND2_X1 _37109_ (.A1(_11954_),
    .A2(_11948_),
    .ZN(_18642_));
 AND2_X1 _37110_ (.A1(_11851_),
    .A2(_11953_),
    .ZN(_18643_));
 AND2_X1 _37111_ (.A1(_11852_),
    .A2(_11951_),
    .ZN(_18641_));
 AND2_X1 _37112_ (.A1(_11651_),
    .A2(_11879_),
    .ZN(_17657_));
 NOR2_X1 _37113_ (.A1(_15196_),
    .A2(_18712_),
    .ZN(_17658_));
 AND2_X1 _37114_ (.A1(_11645_),
    .A2(_11881_),
    .ZN(_17667_));
 AND2_X1 _37115_ (.A1(_11888_),
    .A2(_11886_),
    .ZN(_17666_));
 AND2_X1 _37116_ (.A1(_11648_),
    .A2(_11878_),
    .ZN(_17661_));
 AND2_X1 _37117_ (.A1(_11651_),
    .A2(_11880_),
    .ZN(_17662_));
 AND2_X1 _37118_ (.A1(_11654_),
    .A2(_11879_),
    .ZN(_17663_));
 BUF_X2 _37119_ (.A(net353),
    .Z(_11968_));
 INV_X2 _37120_ (.A(_11968_),
    .ZN(_19029_));
 NOR2_X1 _37121_ (.A1(_18850_),
    .A2(_19029_),
    .ZN(_18368_));
 BUF_X2 _37122_ (.A(a[119]),
    .Z(_11969_));
 AND2_X1 _37123_ (.A1(_11916_),
    .A2(_11969_),
    .ZN(_17684_));
 BUF_X2 _37124_ (.A(net19),
    .Z(_11970_));
 AND2_X1 _37125_ (.A1(_11926_),
    .A2(_11970_),
    .ZN(_17683_));
 INV_X2 _37126_ (.A(_11969_),
    .ZN(_17670_));
 NOR2_X1 _37127_ (.A1(_18850_),
    .A2(_17670_),
    .ZN(_17681_));
 BUF_X2 _37128_ (.A(net21),
    .Z(_11971_));
 AND2_X1 _37129_ (.A1(_11678_),
    .A2(_11971_),
    .ZN(_18257_));
 NOR2_X1 _37130_ (.A1(_14944_),
    .A2(_19029_),
    .ZN(_18258_));
 AND2_X1 _37131_ (.A1(_11916_),
    .A2(_11970_),
    .ZN(_18267_));
 BUF_X2 _37132_ (.A(net18),
    .Z(_11972_));
 AND2_X1 _37133_ (.A1(_11926_),
    .A2(_11972_),
    .ZN(_18266_));
 AND2_X1 _37134_ (.A1(_11928_),
    .A2(_11968_),
    .ZN(_18261_));
 AND2_X1 _37135_ (.A1(_11678_),
    .A2(_11969_),
    .ZN(_18262_));
 AND2_X1 _37136_ (.A1(_11929_),
    .A2(_11971_),
    .ZN(_18263_));
 AND2_X1 _37137_ (.A1(_11670_),
    .A2(_11972_),
    .ZN(_17687_));
 AND2_X1 _37138_ (.A1(_11926_),
    .A2(_11961_),
    .ZN(_17688_));
 AND2_X1 _37139_ (.A1(_11670_),
    .A2(_11961_),
    .ZN(_17708_));
 AND2_X1 _37140_ (.A1(_11926_),
    .A2(_11962_),
    .ZN(_17709_));
 AND2_X1 _37141_ (.A1(_11928_),
    .A2(_11971_),
    .ZN(_17695_));
 AND2_X1 _37142_ (.A1(_11678_),
    .A2(_11970_),
    .ZN(_17696_));
 NOR2_X1 _37143_ (.A1(_14944_),
    .A2(_17670_),
    .ZN(_17697_));
 AND2_X1 _37144_ (.A1(_11678_),
    .A2(_11961_),
    .ZN(_21005_));
 AND2_X1 _37145_ (.A1(_11929_),
    .A2(_11972_),
    .ZN(_21006_));
 AND2_X1 _37146_ (.A1(_11929_),
    .A2(_11961_),
    .ZN(_21008_));
 AND2_X1 _37147_ (.A1(_11678_),
    .A2(_11962_),
    .ZN(_21007_));
 AND2_X1 _37148_ (.A1(_11670_),
    .A2(_11962_),
    .ZN(_17704_));
 AND2_X1 _37149_ (.A1(_11926_),
    .A2(_11960_),
    .ZN(_17705_));
 AND2_X1 _37150_ (.A1(_11928_),
    .A2(_11970_),
    .ZN(_17745_));
 AND2_X1 _37151_ (.A1(_11925_),
    .A2(_11971_),
    .ZN(_17746_));
 AND2_X1 _37152_ (.A1(_11930_),
    .A2(_11969_),
    .ZN(_17747_));
 AND2_X1 _37153_ (.A1(_11670_),
    .A2(_11960_),
    .ZN(_17737_));
 AND2_X1 _37154_ (.A1(_11926_),
    .A2(_11877_),
    .ZN(_17738_));
 AND2_X1 _37155_ (.A1(_11928_),
    .A2(_11969_),
    .ZN(_17721_));
 AND2_X1 _37156_ (.A1(_11678_),
    .A2(_11972_),
    .ZN(_17720_));
 AND2_X1 _37157_ (.A1(_11929_),
    .A2(_11970_),
    .ZN(_17722_));
 AND2_X1 _37158_ (.A1(_11930_),
    .A2(_11971_),
    .ZN(_17725_));
 NOR2_X1 _37159_ (.A1(_14888_),
    .A2(_19029_),
    .ZN(_17726_));
 AND2_X1 _37160_ (.A1(_11673_),
    .A2(_11876_),
    .ZN(_21009_));
 AND2_X1 _37161_ (.A1(_11670_),
    .A2(_11877_),
    .ZN(_21010_));
 NOR2_X1 _37162_ (.A1(_14888_),
    .A2(_17670_),
    .ZN(_17767_));
 AND2_X1 _37163_ (.A1(_11928_),
    .A2(_11972_),
    .ZN(_17766_));
 AND2_X1 _37164_ (.A1(_11930_),
    .A2(_11970_),
    .ZN(_17768_));
 AND2_X1 _37165_ (.A1(_11927_),
    .A2(_11971_),
    .ZN(_17771_));
 NOR2_X1 _37166_ (.A1(_14841_),
    .A2(_19029_),
    .ZN(_17772_));
 AND2_X1 _37167_ (.A1(_11678_),
    .A2(_11960_),
    .ZN(_17783_));
 AND2_X1 _37168_ (.A1(_11684_),
    .A2(_11961_),
    .ZN(_17784_));
 AND2_X1 _37169_ (.A1(_11929_),
    .A2(_11962_),
    .ZN(_17785_));
 AND2_X1 _37170_ (.A1(_11930_),
    .A2(_11972_),
    .ZN(_17794_));
 AND2_X1 _37171_ (.A1(_11927_),
    .A2(_11969_),
    .ZN(_17793_));
 AND2_X1 _37172_ (.A1(_11925_),
    .A2(_11970_),
    .ZN(_17792_));
 AND2_X1 _37173_ (.A1(_11929_),
    .A2(_11960_),
    .ZN(_18206_));
 AND2_X1 _37174_ (.A1(_11670_),
    .A2(_11876_),
    .ZN(_18205_));
 AND2_X1 _37175_ (.A1(_11678_),
    .A2(_11877_),
    .ZN(_18207_));
 AND2_X1 _37176_ (.A1(_11927_),
    .A2(_11970_),
    .ZN(_21051_));
 NOR2_X1 _37177_ (.A1(_14841_),
    .A2(_17670_),
    .ZN(_21052_));
 AND2_X1 _37178_ (.A1(_11693_),
    .A2(_11972_),
    .ZN(_18211_));
 AND2_X1 _37179_ (.A1(_11684_),
    .A2(_11962_),
    .ZN(_18210_));
 AND2_X1 _37180_ (.A1(_11930_),
    .A2(_11961_),
    .ZN(_18209_));
 AND2_X1 _37181_ (.A1(_11693_),
    .A2(_11961_),
    .ZN(_21012_));
 AND2_X1 _37182_ (.A1(_11930_),
    .A2(_11962_),
    .ZN(_21013_));
 AND2_X1 _37183_ (.A1(_11684_),
    .A2(_11877_),
    .ZN(_21015_));
 AND2_X1 _37184_ (.A1(_11929_),
    .A2(_11876_),
    .ZN(_21016_));
 AND2_X1 _37185_ (.A1(_11684_),
    .A2(_11960_),
    .ZN(_17797_));
 AND2_X1 _37186_ (.A1(_11678_),
    .A2(_11876_),
    .ZN(_17799_));
 AND2_X1 _37187_ (.A1(_11929_),
    .A2(_11877_),
    .ZN(_17798_));
 AND2_X1 _37188_ (.A1(_11781_),
    .A2(_11969_),
    .ZN(_17807_));
 AND2_X1 _37189_ (.A1(_11927_),
    .A2(_11972_),
    .ZN(_17806_));
 AND2_X1 _37190_ (.A1(_11931_),
    .A2(_11970_),
    .ZN(_17808_));
 AND2_X1 _37191_ (.A1(_11691_),
    .A2(_11961_),
    .ZN(_17816_));
 AND2_X1 _37192_ (.A1(_11726_),
    .A2(_11960_),
    .ZN(_17817_));
 AND2_X1 _37193_ (.A1(_11693_),
    .A2(_11962_),
    .ZN(_17818_));
 AND2_X1 _37194_ (.A1(_11691_),
    .A2(_11877_),
    .ZN(_21018_));
 AND2_X1 _37195_ (.A1(_11693_),
    .A2(_11876_),
    .ZN(_21019_));
 AND2_X1 _37196_ (.A1(_11931_),
    .A2(_11960_),
    .ZN(_19034_));
 AND2_X1 _37197_ (.A1(_11781_),
    .A2(_11962_),
    .ZN(_19035_));
 NOR2_X1 _37198_ (.A1(_18805_),
    .A2(_18987_),
    .ZN(_17821_));
 AND2_X1 _37199_ (.A1(_11943_),
    .A2(_11965_),
    .ZN(_18183_));
 AND2_X1 _37200_ (.A1(_11939_),
    .A2(_11964_),
    .ZN(_18184_));
 NOR2_X1 _37201_ (.A1(_18805_),
    .A2(_18314_),
    .ZN(_18180_));
 AND2_X1 _37202_ (.A1(_11941_),
    .A2(_11965_),
    .ZN(_17824_));
 AND2_X1 _37203_ (.A1(_11698_),
    .A2(_11967_),
    .ZN(_17825_));
 AND2_X1 _37204_ (.A1(_11709_),
    .A2(_11963_),
    .ZN(_17826_));
 AND2_X1 _37205_ (.A1(_11943_),
    .A2(_11964_),
    .ZN(_17830_));
 AND2_X1 _37206_ (.A1(_11939_),
    .A2(_11966_),
    .ZN(_17829_));
 AND2_X1 _37207_ (.A1(_11698_),
    .A2(_11963_),
    .ZN(_17848_));
 AND2_X1 _37208_ (.A1(_11706_),
    .A2(_11964_),
    .ZN(_17849_));
 NOR2_X1 _37209_ (.A1(_15651_),
    .A2(_18314_),
    .ZN(_17850_));
 AND2_X1 _37210_ (.A1(_11943_),
    .A2(_11966_),
    .ZN(_17846_));
 AND2_X1 _37211_ (.A1(_11939_),
    .A2(_11957_),
    .ZN(_17845_));
 NOR2_X1 _37212_ (.A1(_14677_),
    .A2(_18314_),
    .ZN(_21023_));
 AND2_X1 _37213_ (.A1(_11947_),
    .A2(_11964_),
    .ZN(_21022_));
 AND2_X1 _37214_ (.A1(_11703_),
    .A2(_11872_),
    .ZN(_17893_));
 AND2_X1 _37215_ (.A1(_11709_),
    .A2(_11958_),
    .ZN(_17894_));
 AND2_X1 _37216_ (.A1(_11706_),
    .A2(_11871_),
    .ZN(_17895_));
 AND2_X1 _37217_ (.A1(_11698_),
    .A2(_11959_),
    .ZN(_17899_));
 AND2_X1 _37218_ (.A1(_11945_),
    .A2(_11966_),
    .ZN(_17898_));
 AND2_X1 _37219_ (.A1(_11701_),
    .A2(_11957_),
    .ZN(_17897_));
 AND2_X1 _37220_ (.A1(_11945_),
    .A2(_11957_),
    .ZN(_21025_));
 AND2_X1 _37221_ (.A1(_11701_),
    .A2(_11959_),
    .ZN(_21026_));
 AND2_X1 _37222_ (.A1(_11698_),
    .A2(_11958_),
    .ZN(_17908_));
 AND2_X1 _37223_ (.A1(_11706_),
    .A2(_11872_),
    .ZN(_17907_));
 AND2_X1 _37224_ (.A1(_11709_),
    .A2(_11871_),
    .ZN(_17906_));
 AND2_X1 _37225_ (.A1(_11947_),
    .A2(_11966_),
    .ZN(_17920_));
 AND2_X1 _37226_ (.A1(_11946_),
    .A2(_11965_),
    .ZN(_17921_));
 AND2_X1 _37227_ (.A1(_11873_),
    .A2(_11964_),
    .ZN(_17922_));
 AND2_X1 _37228_ (.A1(_11709_),
    .A2(_11872_),
    .ZN(_21030_));
 AND2_X1 _37229_ (.A1(_11698_),
    .A2(_11871_),
    .ZN(_21029_));
 AND2_X1 _37230_ (.A1(_11947_),
    .A2(_11957_),
    .ZN(_18159_));
 AND2_X1 _37231_ (.A1(_11701_),
    .A2(_11958_),
    .ZN(_18158_));
 AND2_X1 _37232_ (.A1(_11695_),
    .A2(_11959_),
    .ZN(_18157_));
 AND2_X1 _37233_ (.A1(_11663_),
    .A2(_11685_),
    .ZN(_21032_));
 AND2_X1 _37234_ (.A1(_11893_),
    .A2(_11686_),
    .ZN(_21033_));
 AND2_X1 _37235_ (.A1(_11891_),
    .A2(_11884_),
    .ZN(_18718_));
 AND2_X1 _37236_ (.A1(_11857_),
    .A2(_11883_),
    .ZN(_18719_));
 AND2_X1 _37237_ (.A1(_11701_),
    .A2(_11940_),
    .ZN(_17997_));
 AND2_X1 _37238_ (.A1(_11947_),
    .A2(_11937_),
    .ZN(_17996_));
 AND2_X1 _37239_ (.A1(_11695_),
    .A2(_11938_),
    .ZN(_17995_));
 NOR2_X1 _37240_ (.A1(_18805_),
    .A2(_18804_),
    .ZN(_18533_));
 AND2_X1 _37241_ (.A1(_11726_),
    .A2(_11924_),
    .ZN(_18044_));
 AND2_X1 _37242_ (.A1(_11691_),
    .A2(_11922_),
    .ZN(_18043_));
 AND2_X1 _37243_ (.A1(_11693_),
    .A2(_11923_),
    .ZN(_18042_));
 AND2_X1 _37244_ (.A1(_11857_),
    .A2(_11913_),
    .ZN(_18072_));
 AND2_X1 _37245_ (.A1(_11657_),
    .A2(_11915_),
    .ZN(_18073_));
 AND2_X1 _37246_ (.A1(_11891_),
    .A2(_11914_),
    .ZN(_18074_));
 AND2_X1 _37247_ (.A1(_11663_),
    .A2(_11814_),
    .ZN(_21071_));
 AND2_X1 _37248_ (.A1(_11657_),
    .A2(_11813_),
    .ZN(_21070_));
 AND2_X1 _37249_ (.A1(_11663_),
    .A2(_11909_),
    .ZN(_18111_));
 AND2_X1 _37250_ (.A1(_11648_),
    .A2(_11910_),
    .ZN(_18110_));
 AND2_X1 _37251_ (.A1(_11660_),
    .A2(_11911_),
    .ZN(_18112_));
 AND2_X1 _37252_ (.A1(_11907_),
    .A2(_11903_),
    .ZN(_18122_));
 AND2_X1 _37253_ (.A1(_11809_),
    .A2(_11847_),
    .ZN(_18123_));
 AND2_X1 _37254_ (.A1(_11802_),
    .A2(_11846_),
    .ZN(_18124_));
 AND2_X1 _37255_ (.A1(_11802_),
    .A2(_11847_),
    .ZN(_21076_));
 AND2_X1 _37256_ (.A1(_11907_),
    .A2(_11846_),
    .ZN(_21075_));
 AND2_X1 _37257_ (.A1(_11954_),
    .A2(_11902_),
    .ZN(_21048_));
 AND2_X1 _37258_ (.A1(_11852_),
    .A2(_11901_),
    .ZN(_21049_));
 AND2_X1 _37259_ (.A1(_11851_),
    .A2(_11901_),
    .ZN(_18423_));
 AND2_X1 _37260_ (.A1(_11954_),
    .A2(_11903_),
    .ZN(_18424_));
 AND2_X1 _37261_ (.A1(_11765_),
    .A2(_11902_),
    .ZN(_18425_));
 AND2_X1 _37262_ (.A1(_11698_),
    .A2(_11872_),
    .ZN(_18172_));
 AND2_X1 _37263_ (.A1(_11695_),
    .A2(_11958_),
    .ZN(_18173_));
 AND2_X1 _37264_ (.A1(_11701_),
    .A2(_11871_),
    .ZN(_18171_));
 AND2_X1 _37265_ (.A1(_11873_),
    .A2(_11957_),
    .ZN(_21065_));
 AND2_X1 _37266_ (.A1(_11947_),
    .A2(_11959_),
    .ZN(_21066_));
 AND2_X1 _37267_ (.A1(_11706_),
    .A2(_11963_),
    .ZN(_18192_));
 NOR2_X1 _37268_ (.A1(_15651_),
    .A2(_18987_),
    .ZN(_18193_));
 AND2_X1 _37269_ (.A1(_11660_),
    .A2(_11884_),
    .ZN(_18238_));
 AND2_X1 _37270_ (.A1(_11657_),
    .A2(_11882_),
    .ZN(_18237_));
 AND2_X1 _37271_ (.A1(_11663_),
    .A2(_11883_),
    .ZN(_18236_));
 AND2_X1 _37272_ (.A1(_11695_),
    .A2(_11771_),
    .ZN(_21057_));
 AND2_X1 _37273_ (.A1(_11716_),
    .A2(_11773_),
    .ZN(_21058_));
 AND2_X1 _37274_ (.A1(_11873_),
    .A2(_11940_),
    .ZN(_18810_));
 AND2_X1 _37275_ (.A1(_11946_),
    .A2(_11938_),
    .ZN(_18809_));
 AND2_X1 _37276_ (.A1(_11693_),
    .A2(_11795_),
    .ZN(_21060_));
 AND2_X1 _37277_ (.A1(_11691_),
    .A2(_11794_),
    .ZN(_21059_));
 AND2_X1 _37278_ (.A1(_11931_),
    .A2(_11924_),
    .ZN(_18855_));
 AND2_X1 _37279_ (.A1(_11781_),
    .A2(_11923_),
    .ZN(_18856_));
 NOR2_X1 _37280_ (.A1(_18850_),
    .A2(_18849_),
    .ZN(_18582_));
 AND2_X1 _37281_ (.A1(_11643_),
    .A2(_11911_),
    .ZN(_18250_));
 AND2_X1 _37282_ (.A1(_11645_),
    .A2(_11908_),
    .ZN(_18246_));
 AND2_X1 _37283_ (.A1(_11643_),
    .A2(_11909_),
    .ZN(_18245_));
 NOR2_X1 _37284_ (.A1(_18757_),
    .A2(_18945_),
    .ZN(_18484_));
 AND2_X1 _37285_ (.A1(_11873_),
    .A2(_11958_),
    .ZN(_18992_));
 AND2_X1 _37286_ (.A1(_11946_),
    .A2(_11959_),
    .ZN(_18993_));
 AND2_X1 _37287_ (.A1(_11891_),
    .A2(_11915_),
    .ZN(_18903_));
 AND2_X1 _37288_ (.A1(_11857_),
    .A2(_11914_),
    .ZN(_18904_));
 NOR2_X1 _37289_ (.A1(_18757_),
    .A2(_18756_),
    .ZN(_18686_));
 INV_X1 _37290_ (.A(_19483_),
    .ZN(_14226_));
 INV_X1 _37291_ (.A(_19540_),
    .ZN(_14245_));
 INV_X1 _37292_ (.A(_19654_),
    .ZN(_14283_));
 INV_X1 _37293_ (.A(_19825_),
    .ZN(_14334_));
 INV_X1 _37294_ (.A(_19939_),
    .ZN(_14368_));
 INV_X1 _37295_ (.A(_20224_),
    .ZN(_14453_));
 INV_X1 _37296_ (.A(_20281_),
    .ZN(_14470_));
 INV_X1 _37297_ (.A(_20334_),
    .ZN(_14474_));
 BUF_X4 _37298_ (.A(_11665_),
    .Z(_11973_));
 NAND2_X1 _37299_ (.A1(_11751_),
    .A2(_11973_),
    .ZN(_14522_));
 NAND2_X1 _37300_ (.A1(_11751_),
    .A2(_11668_),
    .ZN(_14560_));
 NAND2_X1 _37301_ (.A1(_11717_),
    .A2(_11777_),
    .ZN(_14695_));
 CLKBUF_X3 _37302_ (.A(_11727_),
    .Z(_11974_));
 NAND2_X1 _37303_ (.A1(_11974_),
    .A2(_11739_),
    .ZN(_14719_));
 BUF_X4 _37304_ (.A(_11688_),
    .Z(_11975_));
 NAND2_X1 _37305_ (.A1(_11975_),
    .A2(_11742_),
    .ZN(_14779_));
 INV_X1 _37306_ (.A(_20703_),
    .ZN(_15033_));
 CLKBUF_X3 _37307_ (.A(_11776_),
    .Z(_11976_));
 NAND2_X1 _37308_ (.A1(_11976_),
    .A2(_11783_),
    .ZN(_15363_));
 NAND2_X1 _37309_ (.A1(_11976_),
    .A2(_11785_),
    .ZN(_15381_));
 INV_X1 _37310_ (.A(_20745_),
    .ZN(_15430_));
 NAND2_X1 _37311_ (.A1(_11681_),
    .A2(_11728_),
    .ZN(_15483_));
 INV_X1 _37312_ (.A(_20772_),
    .ZN(_15718_));
 NAND2_X1 _37313_ (.A1(_11766_),
    .A2(_11816_),
    .ZN(_15731_));
 BUF_X4 _37314_ (.A(_11803_),
    .Z(_11977_));
 NAND2_X1 _37315_ (.A1(_11977_),
    .A2(_11826_),
    .ZN(_15771_));
 NAND2_X1 _37316_ (.A1(_11977_),
    .A2(_11833_),
    .ZN(_16129_));
 NAND2_X1 _37317_ (.A1(_11977_),
    .A2(_11832_),
    .ZN(_16166_));
 NAND2_X1 _37318_ (.A1(_11766_),
    .A2(_11836_),
    .ZN(_16206_));
 NAND2_X1 _37319_ (.A1(_11977_),
    .A2(_11836_),
    .ZN(_16214_));
 INV_X1 _37320_ (.A(_20825_),
    .ZN(_16234_));
 NAND2_X1 _37321_ (.A1(_11973_),
    .A2(_11861_),
    .ZN(_16239_));
 BUF_X4 _37322_ (.A(_11667_),
    .Z(_11978_));
 NAND2_X1 _37323_ (.A1(_11978_),
    .A2(_11868_),
    .ZN(_16285_));
 NAND2_X1 _37324_ (.A1(_11699_),
    .A2(_11777_),
    .ZN(_16547_));
 NAND2_X1 _37325_ (.A1(_11973_),
    .A2(_11879_),
    .ZN(_16652_));
 NAND2_X1 _37326_ (.A1(_11978_),
    .A2(_11879_),
    .ZN(_16671_));
 NAND2_X1 _37327_ (.A1(_11978_),
    .A2(_11886_),
    .ZN(_16685_));
 INV_X1 _37328_ (.A(_20858_),
    .ZN(_16718_));
 NAND2_X1 _37329_ (.A1(_11977_),
    .A2(_11896_),
    .ZN(_16819_));
 NAND2_X1 _37330_ (.A1(_11978_),
    .A2(_11910_),
    .ZN(_16966_));
 NAND2_X1 _37331_ (.A1(_11975_),
    .A2(_11919_),
    .ZN(_17063_));
 NAND2_X1 _37332_ (.A1(_11976_),
    .A2(_11934_),
    .ZN(_17200_));
 INV_X1 _37333_ (.A(_20950_),
    .ZN(_17233_));
 NAND2_X1 _37334_ (.A1(_11976_),
    .A2(_11936_),
    .ZN(_17247_));
 INV_X1 _37335_ (.A(_20959_),
    .ZN(_17289_));
 NAND2_X1 _37336_ (.A1(_11974_),
    .A2(_11972_),
    .ZN(_17436_));
 NAND2_X1 _37337_ (.A1(_11977_),
    .A2(_11952_),
    .ZN(_17635_));
 INV_X1 _37338_ (.A(_21021_),
    .ZN(_17901_));
 INV_X1 _37339_ (.A(_21047_),
    .ZN(_18127_));
 INV_X1 _37340_ (.A(_20981_),
    .ZN(_18277_));
 NAND2_X1 _37341_ (.A1(_11975_),
    .A2(_11972_),
    .ZN(_18327_));
 NAND2_X1 _37342_ (.A1(_11977_),
    .A2(_11950_),
    .ZN(_18649_));
 NAND2_X1 _37343_ (.A1(_11973_),
    .A2(_11649_),
    .ZN(_19076_));
 BUF_X4 _37344_ (.A(_11718_),
    .Z(_11979_));
 NAND2_X1 _37345_ (.A1(_11711_),
    .A2(_11979_),
    .ZN(_19169_));
 NAND2_X1 _37346_ (.A1(_11973_),
    .A2(_11856_),
    .ZN(_19257_));
 NAND2_X1 _37347_ (.A1(_11766_),
    .A2(_11806_),
    .ZN(_19307_));
 NAND2_X1 _37348_ (.A1(_11979_),
    .A2(_11779_),
    .ZN(_19357_));
 NAND2_X1 _37349_ (.A1(_11733_),
    .A2(_11728_),
    .ZN(_19401_));
 INV_X1 _37350_ (.A(_19882_),
    .ZN(_14351_));
 INV_X1 _37351_ (.A(_20648_),
    .ZN(_14561_));
 NAND2_X1 _37352_ (.A1(_11679_),
    .A2(_11671_),
    .ZN(_14570_));
 NAND2_X1 _37353_ (.A1(_11973_),
    .A2(_11658_),
    .ZN(_14617_));
 NAND2_X1 _37354_ (.A1(_11978_),
    .A2(_11658_),
    .ZN(_14629_));
 NAND2_X1 _37355_ (.A1(_11974_),
    .A2(_11738_),
    .ZN(_14715_));
 NAND2_X1 _37356_ (.A1(_11975_),
    .A2(_11738_),
    .ZN(_14720_));
 NAND2_X1 _37357_ (.A1(_11974_),
    .A2(_11742_),
    .ZN(_14766_));
 NAND2_X1 _37358_ (.A1(_11730_),
    .A2(_11743_),
    .ZN(_14842_));
 NAND2_X1 _37359_ (.A1(_11671_),
    .A2(_11743_),
    .ZN(_14958_));
 NAND2_X1 _37360_ (.A1(_11676_),
    .A2(_11975_),
    .ZN(_15020_));
 NAND2_X1 _37361_ (.A1(_11676_),
    .A2(_11728_),
    .ZN(_15034_));
 NAND2_X1 _37362_ (.A1(_11749_),
    .A2(_11752_),
    .ZN(_15156_));
 NAND2_X1 _37363_ (.A1(_11679_),
    .A2(_11740_),
    .ZN(_15176_));
 NAND2_X1 _37364_ (.A1(_11752_),
    .A2(_11748_),
    .ZN(_15197_));
 NAND2_X1 _37365_ (.A1(_11752_),
    .A2(_11747_),
    .ZN(_15239_));
 NAND2_X1 _37366_ (.A1(_11752_),
    .A2(_11664_),
    .ZN(_15314_));
 NAND2_X1 _37367_ (.A1(_11724_),
    .A2(_11717_),
    .ZN(_15413_));
 NAND2_X1 _37368_ (.A1(_11976_),
    .A2(_11788_),
    .ZN(_15431_));
 NAND2_X1 _37369_ (.A1(_11979_),
    .A2(_11788_),
    .ZN(_15460_));
 INV_X1 _37370_ (.A(_20738_),
    .ZN(_15484_));
 NAND2_X1 _37371_ (.A1(_11681_),
    .A2(_11975_),
    .ZN(_15604_));
 NAND2_X1 _37372_ (.A1(_11977_),
    .A2(_11816_),
    .ZN(_15719_));
 INV_X1 _37373_ (.A(_20780_),
    .ZN(_15772_));
 NAND2_X1 _37374_ (.A1(_11766_),
    .A2(_11826_),
    .ZN(_15807_));
 NAND2_X1 _37375_ (.A1(_11823_),
    .A2(_11827_),
    .ZN(_15916_));
 NAND2_X1 _37376_ (.A1(_11830_),
    .A2(_11827_),
    .ZN(_15965_));
 INV_X1 _37377_ (.A(_20803_),
    .ZN(_16167_));
 NAND2_X1 _37378_ (.A1(_11978_),
    .A2(_11863_),
    .ZN(_16240_));
 INV_X1 _37379_ (.A(_20833_),
    .ZN(_16286_));
 NAND2_X1 _37380_ (.A1(_11973_),
    .A2(_11868_),
    .ZN(_16295_));
 NAND2_X1 _37381_ (.A1(_11664_),
    .A2(_11869_),
    .ZN(_16362_));
 NAND2_X1 _37382_ (.A1(_11720_),
    .A2(_11717_),
    .ZN(_16473_));
 NAND2_X1 _37383_ (.A1(_11749_),
    .A2(_11869_),
    .ZN(_16486_));
 NAND2_X1 _37384_ (.A1(_11696_),
    .A2(_11777_),
    .ZN(_16556_));
 NAND2_X1 _37385_ (.A1(_11747_),
    .A2(_11878_),
    .ZN(_16601_));
 INV_X1 _37386_ (.A(_20875_),
    .ZN(_16672_));
 NAND2_X1 _37387_ (.A1(_11714_),
    .A2(_11777_),
    .ZN(_16719_));
 NAND2_X1 _37388_ (.A1(_11713_),
    .A2(_11714_),
    .ZN(_16723_));
 NAND2_X1 _37389_ (.A1(_11823_),
    .A2(_11895_),
    .ZN(_16786_));
 NAND2_X1 _37390_ (.A1(_11763_),
    .A2(_11895_),
    .ZN(_16816_));
 INV_X1 _37391_ (.A(_20897_),
    .ZN(_16820_));
 NAND2_X1 _37392_ (.A1(_11973_),
    .A2(_11909_),
    .ZN(_16905_));
 NAND2_X1 _37393_ (.A1(_11973_),
    .A2(_11912_),
    .ZN(_16967_));
 NAND2_X1 _37394_ (.A1(_11674_),
    .A2(_11919_),
    .ZN(_16976_));
 NAND2_X1 _37395_ (.A1(_11740_),
    .A2(_11920_),
    .ZN(_17025_));
 INV_X1 _37396_ (.A(_20931_),
    .ZN(_17096_));
 NAND2_X1 _37397_ (.A1(_11974_),
    .A2(_11921_),
    .ZN(_17110_));
 NAND2_X1 _37398_ (.A1(_11979_),
    .A2(_11935_),
    .ZN(_17201_));
 NAND2_X1 _37399_ (.A1(_11976_),
    .A2(_11935_),
    .ZN(_17234_));
 NAND2_X1 _37400_ (.A1(_11977_),
    .A2(_11956_),
    .ZN(_17276_));
 NAND2_X1 _37401_ (.A1(_11977_),
    .A2(_11955_),
    .ZN(_17290_));
 NAND2_X1 _37402_ (.A1(_11763_),
    .A2(_11956_),
    .ZN(_17337_));
 NAND2_X1 _37403_ (.A1(_11837_),
    .A2(_11955_),
    .ZN(_17349_));
 NAND2_X1 _37404_ (.A1(_11766_),
    .A2(_11896_),
    .ZN(_17544_));
 INV_X1 _37405_ (.A(_20917_),
    .ZN(_17553_));
 NAND2_X1 _37406_ (.A1(_11748_),
    .A2(_11878_),
    .ZN(_17653_));
 NAND2_X1 _37407_ (.A1(_11671_),
    .A2(_11968_),
    .ZN(_17671_));
 NAND2_X1 _37408_ (.A1(_11740_),
    .A2(_11968_),
    .ZN(_17691_));
 NAND2_X1 _37409_ (.A1(_11975_),
    .A2(_11971_),
    .ZN(_17789_));
 NAND2_X1 _37410_ (.A1(_11724_),
    .A2(_11967_),
    .ZN(_17842_));
 NAND2_X1 _37411_ (.A1(_11979_),
    .A2(_11963_),
    .ZN(_17867_));
 NAND2_X1 _37412_ (.A1(_11976_),
    .A2(_11963_),
    .ZN(_17902_));
 NAND2_X1 _37413_ (.A1(_11804_),
    .A2(_11900_),
    .ZN(_18128_));
 NAND2_X1 _37414_ (.A1(_11979_),
    .A2(_11966_),
    .ZN(_18167_));
 NAND2_X1 _37415_ (.A1(_11720_),
    .A2(_11967_),
    .ZN(_18175_));
 INV_X1 _37416_ (.A(_21014_),
    .ZN(_18219_));
 NAND2_X1 _37417_ (.A1(_11713_),
    .A2(_11963_),
    .ZN(_18315_));
 NAND2_X1 _37418_ (.A1(_11682_),
    .A2(_11968_),
    .ZN(_18361_));
 NAND2_X1 _37419_ (.A1(_11978_),
    .A2(_11912_),
    .ZN(_18372_));
 NAND2_X1 _37420_ (.A1(_11748_),
    .A2(_11908_),
    .ZN(_18416_));
 NAND2_X1 _37421_ (.A1(_11766_),
    .A2(_11900_),
    .ZN(_18437_));
 NAND2_X1 _37422_ (.A1(_11830_),
    .A2(_11895_),
    .ZN(_18481_));
 NAND2_X1 _37423_ (.A1(_11979_),
    .A2(_11936_),
    .ZN(_18493_));
 NAND2_X1 _37424_ (.A1(_11975_),
    .A2(_11921_),
    .ZN(_18542_));
 NAND2_X1 _37425_ (.A1(_11973_),
    .A2(_11886_),
    .ZN(_18594_));
 NAND2_X1 _37426_ (.A1(_11766_),
    .A2(_11952_),
    .ZN(_18650_));
 NAND2_X1 _37427_ (.A1(_11704_),
    .A2(_11777_),
    .ZN(_19170_));
 NAND2_X1 _37428_ (.A1(_11975_),
    .A2(_11753_),
    .ZN(_19214_));
 NAND2_X1 _37429_ (.A1(_11976_),
    .A2(_11780_),
    .ZN(_19358_));
 INV_X1 _37430_ (.A(_19479_),
    .ZN(_14213_));
 INV_X1 _37431_ (.A(_19536_),
    .ZN(_14232_));
 INV_X1 _37432_ (.A(_19593_),
    .ZN(_14251_));
 INV_X1 _37433_ (.A(_19597_),
    .ZN(_14265_));
 INV_X1 _37434_ (.A(_19650_),
    .ZN(_14270_));
 INV_X1 _37435_ (.A(_19707_),
    .ZN(_14289_));
 INV_X1 _37436_ (.A(_19711_),
    .ZN(_14301_));
 INV_X1 _37437_ (.A(_19764_),
    .ZN(_14306_));
 INV_X1 _37438_ (.A(_19768_),
    .ZN(_14318_));
 INV_X1 _37439_ (.A(_19821_),
    .ZN(_14323_));
 INV_X1 _37440_ (.A(_19878_),
    .ZN(_14340_));
 INV_X1 _37441_ (.A(_19935_),
    .ZN(_14357_));
 INV_X1 _37442_ (.A(_19992_),
    .ZN(_14374_));
 INV_X1 _37443_ (.A(_19996_),
    .ZN(_14386_));
 INV_X1 _37444_ (.A(_20049_),
    .ZN(_14391_));
 INV_X1 _37445_ (.A(_20053_),
    .ZN(_14403_));
 INV_X1 _37446_ (.A(_20106_),
    .ZN(_14408_));
 INV_X1 _37447_ (.A(_20110_),
    .ZN(_14420_));
 INV_X1 _37448_ (.A(_20163_),
    .ZN(_14425_));
 INV_X1 _37449_ (.A(_20167_),
    .ZN(_14437_));
 INV_X1 _37450_ (.A(_20220_),
    .ZN(_14442_));
 INV_X1 _37451_ (.A(_20277_),
    .ZN(_14459_));
 INV_X1 _37452_ (.A(_20338_),
    .ZN(_14488_));
 NAND2_X1 _37453_ (.A1(_11752_),
    .A2(_11668_),
    .ZN(_14524_));
 NAND2_X1 _37454_ (.A1(_11676_),
    .A2(_11674_),
    .ZN(_14571_));
 NAND2_X1 _37455_ (.A1(_11978_),
    .A2(_11661_),
    .ZN(_14618_));
 INV_X1 _37456_ (.A(_20660_),
    .ZN(_14630_));
 NAND2_X1 _37457_ (.A1(_11770_),
    .A2(_11717_),
    .ZN(_14679_));
 NAND2_X1 _37458_ (.A1(_11714_),
    .A2(_11979_),
    .ZN(_14697_));
 INV_X1 _37459_ (.A(_20680_),
    .ZN(_14716_));
 INV_X1 _37460_ (.A(_20688_),
    .ZN(_14767_));
 NAND2_X1 _37461_ (.A1(_11974_),
    .A2(_11743_),
    .ZN(_14781_));
 NAND2_X1 _37462_ (.A1(_11740_),
    .A2(_11743_),
    .ZN(_14890_));
 NAND2_X1 _37463_ (.A1(_11682_),
    .A2(_11743_),
    .ZN(_14946_));
 NAND2_X1 _37464_ (.A1(_11674_),
    .A2(_11742_),
    .ZN(_14959_));
 NAND2_X1 _37465_ (.A1(_11679_),
    .A2(_11728_),
    .ZN(_15021_));
 NAND2_X1 _37466_ (.A1(_11679_),
    .A2(_11730_),
    .ZN(_15091_));
 NAND2_X1 _37467_ (.A1(_11751_),
    .A2(_11750_),
    .ZN(_15157_));
 NAND2_X1 _37468_ (.A1(_11679_),
    .A2(_11682_),
    .ZN(_15347_));
 INV_X1 _37469_ (.A(_20732_),
    .ZN(_15365_));
 NAND2_X1 _37470_ (.A1(_11979_),
    .A2(_11783_),
    .ZN(_15383_));
 NAND2_X1 _37471_ (.A1(_11976_),
    .A2(_11789_),
    .ZN(_15461_));
 NAND2_X1 _37472_ (.A1(_11770_),
    .A2(_11789_),
    .ZN(_15537_));
 NAND2_X1 _37473_ (.A1(_11724_),
    .A2(_11789_),
    .ZN(_15579_));
 NAND2_X1 _37474_ (.A1(_11675_),
    .A2(_11728_),
    .ZN(_15605_));
 NAND2_X1 _37475_ (.A1(_11720_),
    .A2(_11789_),
    .ZN(_15653_));
 NAND2_X1 _37476_ (.A1(_11804_),
    .A2(_11818_),
    .ZN(_15733_));
 NAND2_X1 _37477_ (.A1(_11804_),
    .A2(_11827_),
    .ZN(_15808_));
 NAND2_X1 _37478_ (.A1(_11763_),
    .A2(_11827_),
    .ZN(_15872_));
 NAND2_X1 _37479_ (.A1(_11823_),
    .A2(_11833_),
    .ZN(_16026_));
 NAND2_X1 _37480_ (.A1(_11763_),
    .A2(_11833_),
    .ZN(_16086_));
 NAND2_X1 _37481_ (.A1(_11766_),
    .A2(_11832_),
    .ZN(_16131_));
 NAND2_X1 _37482_ (.A1(_11804_),
    .A2(_11834_),
    .ZN(_16208_));
 INV_X1 _37483_ (.A(_20812_),
    .ZN(_16216_));
 NAND2_X1 _37484_ (.A1(_11978_),
    .A2(_11861_),
    .ZN(_16236_));
 NAND2_X1 _37485_ (.A1(_11978_),
    .A2(_11869_),
    .ZN(_16296_));
 NAND2_X1 _37486_ (.A1(_11747_),
    .A2(_11869_),
    .ZN(_16410_));
 NAND2_X1 _37487_ (.A1(_11748_),
    .A2(_11869_),
    .ZN(_16462_));
 NAND2_X1 _37488_ (.A1(_11750_),
    .A2(_11868_),
    .ZN(_16487_));
 NAND2_X1 _37489_ (.A1(_11830_),
    .A2(_11833_),
    .ZN(_16515_));
 NAND2_X1 _37490_ (.A1(_11696_),
    .A2(_11979_),
    .ZN(_16549_));
 INV_X1 _37491_ (.A(_20860_),
    .ZN(_16557_));
 NAND2_X1 _37492_ (.A1(_11664_),
    .A2(_11878_),
    .ZN(_16632_));
 NAND2_X1 _37493_ (.A1(_11668_),
    .A2(_11878_),
    .ZN(_16654_));
 INV_X1 _37494_ (.A(_20884_),
    .ZN(_16687_));
 NAND2_X1 _37495_ (.A1(_11710_),
    .A2(_11717_),
    .ZN(_16724_));
 NAND2_X1 _37496_ (.A1(_11747_),
    .A2(_11908_),
    .ZN(_16889_));
 NAND2_X1 _37497_ (.A1(_11668_),
    .A2(_11908_),
    .ZN(_16906_));
 NAND2_X1 _37498_ (.A1(_11671_),
    .A2(_11920_),
    .ZN(_16977_));
 NAND2_X1 _37499_ (.A1(_11730_),
    .A2(_11920_),
    .ZN(_17056_));
 NAND2_X1 _37500_ (.A1(_11974_),
    .A2(_11920_),
    .ZN(_17065_));
 NAND2_X1 _37501_ (.A1(_11974_),
    .A2(_11919_),
    .ZN(_17097_));
 INV_X1 _37502_ (.A(_20939_),
    .ZN(_17111_));
 NAND2_X1 _37503_ (.A1(_11724_),
    .A2(_11934_),
    .ZN(_17130_));
 NAND2_X1 _37504_ (.A1(_11770_),
    .A2(_11934_),
    .ZN(_17193_));
 INV_X1 _37505_ (.A(_20958_),
    .ZN(_17249_));
 NAND2_X1 _37506_ (.A1(_11766_),
    .A2(_11955_),
    .ZN(_17277_));
 NAND2_X1 _37507_ (.A1(_11831_),
    .A2(_11956_),
    .ZN(_17350_));
 NAND2_X1 _37508_ (.A1(_11823_),
    .A2(_11956_),
    .ZN(_17419_));
 INV_X1 _37509_ (.A(_20982_),
    .ZN(_17438_));
 NAND2_X1 _37510_ (.A1(_11770_),
    .A2(_11967_),
    .ZN(_17464_));
 NAND2_X1 _37511_ (.A1(_11804_),
    .A2(_11895_),
    .ZN(_17545_));
 NAND2_X1 _37512_ (.A1(_11668_),
    .A2(_11909_),
    .ZN(_17554_));
 INV_X1 _37513_ (.A(_21000_),
    .ZN(_17637_));
 NAND2_X1 _37514_ (.A1(_11674_),
    .A2(_11971_),
    .ZN(_17672_));
 NAND2_X1 _37515_ (.A1(_11730_),
    .A2(_11968_),
    .ZN(_17751_));
 NAND2_X1 _37516_ (.A1(_11974_),
    .A2(_11968_),
    .ZN(_17790_));
 NAND2_X1 _37517_ (.A1(_11976_),
    .A2(_11967_),
    .ZN(_17868_));
 NAND2_X1 _37518_ (.A1(_11664_),
    .A2(_11908_),
    .ZN(_18120_));
 NAND2_X1 _37519_ (.A1(_11777_),
    .A2(_11964_),
    .ZN(_18168_));
 NAND2_X1 _37520_ (.A1(_11974_),
    .A2(_11971_),
    .ZN(_18220_));
 NAND2_X1 _37521_ (.A1(_11777_),
    .A2(_11966_),
    .ZN(_18279_));
 NAND2_X1 _37522_ (.A1(_11710_),
    .A2(_11967_),
    .ZN(_18316_));
 NAND2_X1 _37523_ (.A1(_11728_),
    .A2(_11970_),
    .ZN(_18329_));
 INV_X1 _37524_ (.A(_21043_),
    .ZN(_18373_));
 NAND2_X1 _37525_ (.A1(_11804_),
    .A2(_11899_),
    .ZN(_18438_));
 NAND2_X1 _37526_ (.A1(_11777_),
    .A2(_11933_),
    .ZN(_18494_));
 NAND2_X1 _37527_ (.A1(_11720_),
    .A2(_11934_),
    .ZN(_18530_));
 NAND2_X1 _37528_ (.A1(_11728_),
    .A2(_11918_),
    .ZN(_18543_));
 NAND2_X1 _37529_ (.A1(_11682_),
    .A2(_11920_),
    .ZN(_18576_));
 NAND2_X1 _37530_ (.A1(_11668_),
    .A2(_11881_),
    .ZN(_18595_));
 NAND2_X1 _37531_ (.A1(_11830_),
    .A2(_11956_),
    .ZN(_18680_));
 NAND2_X1 _37532_ (.A1(_11668_),
    .A2(_11652_),
    .ZN(_19078_));
 NAND2_X1 _37533_ (.A1(_11728_),
    .A2(_11757_),
    .ZN(_19215_));
 NAND2_X1 _37534_ (.A1(_11668_),
    .A2(_11859_),
    .ZN(_19259_));
 NAND2_X1 _37535_ (.A1(_11807_),
    .A2(_11804_),
    .ZN(_19309_));
 NAND2_X1 _37536_ (.A1(_11975_),
    .A2(_11731_),
    .ZN(_19403_));
 INV_X1 _37537_ (.A(_14531_),
    .ZN(_14537_));
 INV_X1 _37538_ (.A(_14536_),
    .ZN(_14538_));
 INV_X1 _37539_ (.A(_14550_),
    .ZN(_14587_));
 INV_X1 _37540_ (.A(_14555_),
    .ZN(_14588_));
 INV_X1 _37541_ (.A(_14573_),
    .ZN(_19204_));
 INV_X1 _37542_ (.A(_14577_),
    .ZN(_19205_));
 INV_X1 _37543_ (.A(_14581_),
    .ZN(_15350_));
 INV_X1 _37544_ (.A(_14585_),
    .ZN(_15317_));
 INV_X1 _37545_ (.A(_14598_),
    .ZN(_14603_));
 INV_X1 _37546_ (.A(_14602_),
    .ZN(_19091_));
 INV_X1 _37547_ (.A(_14623_),
    .ZN(_19088_));
 INV_X1 _37548_ (.A(_14627_),
    .ZN(_14628_));
 INV_X1 _37549_ (.A(_14641_),
    .ZN(_14654_));
 INV_X1 _37550_ (.A(_14651_),
    .ZN(_16694_));
 INV_X1 _37551_ (.A(_14659_),
    .ZN(_16695_));
 INV_X1 _37552_ (.A(_14668_),
    .ZN(_14682_));
 INV_X1 _37553_ (.A(_14676_),
    .ZN(_14683_));
 INV_X1 _37554_ (.A(_14694_),
    .ZN(_16715_));
 INV_X1 _37555_ (.A(_14703_),
    .ZN(_16716_));
 INV_X1 _37556_ (.A(_14713_),
    .ZN(_14714_));
 INV_X1 _37557_ (.A(_14731_),
    .ZN(_19413_));
 INV_X1 _37558_ (.A(_14740_),
    .ZN(_19416_));
 INV_X1 _37559_ (.A(_14745_),
    .ZN(_14746_));
 INV_X1 _37560_ (.A(_14754_),
    .ZN(_14761_));
 INV_X1 _37561_ (.A(_14759_),
    .ZN(_14762_));
 INV_X1 _37562_ (.A(_14778_),
    .ZN(_14789_));
 INV_X1 _37563_ (.A(_14788_),
    .ZN(_14790_));
 INV_X1 _37564_ (.A(_14795_),
    .ZN(_14796_));
 INV_X1 _37565_ (.A(_14806_),
    .ZN(_14816_));
 INV_X1 _37566_ (.A(_14811_),
    .ZN(_14818_));
 INV_X1 _37567_ (.A(_14815_),
    .ZN(_14817_));
 INV_X1 _37568_ (.A(_14835_),
    .ZN(_14847_));
 INV_X1 _37569_ (.A(_14840_),
    .ZN(_14846_));
 INV_X1 _37570_ (.A(_14861_),
    .ZN(_14873_));
 INV_X1 _37571_ (.A(_14868_),
    .ZN(_14874_));
 INV_X1 _37572_ (.A(_14872_),
    .ZN(_14875_));
 INV_X1 _37573_ (.A(_14887_),
    .ZN(_14898_));
 INV_X1 _37574_ (.A(_14897_),
    .ZN(_14899_));
 INV_X1 _37575_ (.A(_14913_),
    .ZN(_14918_));
 INV_X1 _37576_ (.A(_14917_),
    .ZN(_14919_));
 INV_X1 _37577_ (.A(_14923_),
    .ZN(_14924_));
 INV_X1 _37578_ (.A(_14930_),
    .ZN(_14932_));
 INV_X1 _37579_ (.A(_14939_),
    .ZN(_14940_));
 INV_X1 _37580_ (.A(_14952_),
    .ZN(_14953_));
 INV_X1 _37581_ (.A(_14961_),
    .ZN(_19392_));
 INV_X1 _37582_ (.A(_14964_),
    .ZN(_19393_));
 INV_X1 _37583_ (.A(_14972_),
    .ZN(_14985_));
 INV_X1 _37584_ (.A(_14980_),
    .ZN(_14986_));
 INV_X1 _37585_ (.A(_14984_),
    .ZN(_14987_));
 INV_X1 _37586_ (.A(_15000_),
    .ZN(_15009_));
 INV_X1 _37587_ (.A(_15004_),
    .ZN(_15684_));
 INV_X1 _37588_ (.A(_15008_),
    .ZN(_15685_));
 INV_X1 _37589_ (.A(_15018_),
    .ZN(_15029_));
 INV_X1 _37590_ (.A(_15028_),
    .ZN(_15030_));
 INV_X1 _37591_ (.A(_15041_),
    .ZN(_15672_));
 INV_X1 _37592_ (.A(_15053_),
    .ZN(_15068_));
 INV_X1 _37593_ (.A(_15057_),
    .ZN(_15060_));
 INV_X1 _37594_ (.A(_15066_),
    .ZN(_15067_));
 INV_X1 _37595_ (.A(_15084_),
    .ZN(_15094_));
 INV_X1 _37596_ (.A(_15089_),
    .ZN(_15095_));
 INV_X1 _37597_ (.A(_15110_),
    .ZN(_15120_));
 INV_X1 _37598_ (.A(_15115_),
    .ZN(_15121_));
 INV_X1 _37599_ (.A(_15119_),
    .ZN(_15122_));
 INV_X1 _37600_ (.A(_15138_),
    .ZN(_15150_));
 INV_X1 _37601_ (.A(_15145_),
    .ZN(_15152_));
 INV_X1 _37602_ (.A(_15149_),
    .ZN(_15151_));
 INV_X1 _37603_ (.A(_15159_),
    .ZN(_19067_));
 INV_X1 _37604_ (.A(_15163_),
    .ZN(_19068_));
 INV_X1 _37605_ (.A(_15167_),
    .ZN(_15200_));
 INV_X1 _37606_ (.A(_15171_),
    .ZN(_15218_));
 INV_X1 _37607_ (.A(_15175_),
    .ZN(_15185_));
 INV_X1 _37608_ (.A(_15184_),
    .ZN(_15186_));
 INV_X1 _37609_ (.A(_15208_),
    .ZN(_15222_));
 INV_X1 _37610_ (.A(_15213_),
    .ZN(_15265_));
 INV_X1 _37611_ (.A(_15217_),
    .ZN(_15266_));
 INV_X1 _37612_ (.A(_15234_),
    .ZN(_15269_));
 INV_X1 _37613_ (.A(_15237_),
    .ZN(_15293_));
 INV_X1 _37614_ (.A(_15246_),
    .ZN(_15294_));
 INV_X1 _37615_ (.A(_15251_),
    .ZN(_15256_));
 INV_X1 _37616_ (.A(_15255_),
    .ZN(_15257_));
 INV_X1 _37617_ (.A(_15261_),
    .ZN(_15262_));
 INV_X1 _37618_ (.A(_15280_),
    .ZN(_15309_));
 INV_X1 _37619_ (.A(_15285_),
    .ZN(_15331_));
 INV_X1 _37620_ (.A(_15288_),
    .ZN(_15330_));
 INV_X1 _37621_ (.A(_15292_),
    .ZN(_15332_));
 INV_X1 _37622_ (.A(_15308_),
    .ZN(_15342_));
 INV_X1 _37623_ (.A(_15325_),
    .ZN(_15327_));
 INV_X1 _37624_ (.A(_15362_),
    .ZN(_15364_));
 INV_X1 _37625_ (.A(_15380_),
    .ZN(_19368_));
 INV_X1 _37626_ (.A(_15390_),
    .ZN(_15392_));
 INV_X1 _37627_ (.A(_15399_),
    .ZN(_15402_));
 INV_X1 _37628_ (.A(_15420_),
    .ZN(_15426_));
 INV_X1 _37629_ (.A(_15425_),
    .ZN(_15427_));
 INV_X1 _37630_ (.A(_15442_),
    .ZN(_15449_));
 INV_X1 _37631_ (.A(_15447_),
    .ZN(_15450_));
 INV_X1 _37632_ (.A(_15455_),
    .ZN(_15456_));
 INV_X1 _37633_ (.A(_15468_),
    .ZN(_15475_));
 INV_X1 _37634_ (.A(_15473_),
    .ZN(_15474_));
 INV_X1 _37635_ (.A(_15482_),
    .ZN(_15485_));
 INV_X1 _37636_ (.A(_15499_),
    .ZN(_15513_));
 INV_X1 _37637_ (.A(_15503_),
    .ZN(_15506_));
 INV_X1 _37638_ (.A(_15512_),
    .ZN(_15514_));
 INV_X1 _37639_ (.A(_15527_),
    .ZN(_15540_));
 INV_X1 _37640_ (.A(_15535_),
    .ZN(_15541_));
 INV_X1 _37641_ (.A(_15554_),
    .ZN(_15567_));
 INV_X1 _37642_ (.A(_15561_),
    .ZN(_15568_));
 INV_X1 _37643_ (.A(_15565_),
    .ZN(_15566_));
 INV_X1 _37644_ (.A(_15585_),
    .ZN(_15592_));
 INV_X1 _37645_ (.A(_15590_),
    .ZN(_15591_));
 INV_X1 _37646_ (.A(_15602_),
    .ZN(_19224_));
 INV_X1 _37647_ (.A(_15609_),
    .ZN(_15610_));
 INV_X1 _37648_ (.A(_15617_),
    .ZN(_15622_));
 INV_X1 _37649_ (.A(_15621_),
    .ZN(_15623_));
 INV_X1 _37650_ (.A(_15629_),
    .ZN(_15630_));
 INV_X1 _37651_ (.A(_15637_),
    .ZN(_15638_));
 INV_X1 _37652_ (.A(_15646_),
    .ZN(_15648_));
 INV_X1 _37653_ (.A(_15658_),
    .ZN(_19344_));
 INV_X1 _37654_ (.A(_15662_),
    .ZN(_19345_));
 INV_X1 _37655_ (.A(_15667_),
    .ZN(_15669_));
 INV_X1 _37656_ (.A(_15679_),
    .ZN(_19349_));
 INV_X1 _37657_ (.A(_15691_),
    .ZN(_15697_));
 INV_X1 _37658_ (.A(_15695_),
    .ZN(_15696_));
 INV_X1 _37659_ (.A(_15701_),
    .ZN(_15702_));
 INV_X1 _37660_ (.A(_15717_),
    .ZN(_15720_));
 INV_X1 _37661_ (.A(_15730_),
    .ZN(_19319_));
 INV_X1 _37662_ (.A(_15740_),
    .ZN(_15742_));
 INV_X1 _37663_ (.A(_15753_),
    .ZN(_19322_));
 INV_X1 _37664_ (.A(_15757_),
    .ZN(_15759_));
 INV_X1 _37665_ (.A(_15766_),
    .ZN(_15768_));
 INV_X1 _37666_ (.A(_15784_),
    .ZN(_15791_));
 INV_X1 _37667_ (.A(_15789_),
    .ZN(_15790_));
 INV_X1 _37668_ (.A(_15797_),
    .ZN(_15798_));
 INV_X1 _37669_ (.A(_15805_),
    .ZN(_15816_));
 INV_X1 _37670_ (.A(_15815_),
    .ZN(_15817_));
 INV_X1 _37671_ (.A(_15834_),
    .ZN(_15844_));
 INV_X1 _37672_ (.A(_15839_),
    .ZN(_15845_));
 INV_X1 _37673_ (.A(_15843_),
    .ZN(_15846_));
 INV_X1 _37674_ (.A(_15860_),
    .ZN(_15875_));
 INV_X1 _37675_ (.A(_15864_),
    .ZN(_15867_));
 INV_X1 _37676_ (.A(_15889_),
    .ZN(_15900_));
 INV_X1 _37677_ (.A(_15894_),
    .ZN(_15899_));
 INV_X1 _37678_ (.A(_15898_),
    .ZN(_15901_));
 INV_X1 _37679_ (.A(_15914_),
    .ZN(_15925_));
 INV_X1 _37680_ (.A(_15924_),
    .ZN(_15926_));
 INV_X1 _37681_ (.A(_15933_),
    .ZN(_15938_));
 INV_X1 _37682_ (.A(_15937_),
    .ZN(_15939_));
 INV_X1 _37683_ (.A(_15943_),
    .ZN(_15944_));
 INV_X1 _37684_ (.A(_15950_),
    .ZN(_15953_));
 INV_X1 _37685_ (.A(_15959_),
    .ZN(_15960_));
 INV_X1 _37686_ (.A(_15972_),
    .ZN(_15973_));
 INV_X1 _37687_ (.A(_15979_),
    .ZN(_19294_));
 INV_X1 _37688_ (.A(_15983_),
    .ZN(_19295_));
 INV_X1 _37689_ (.A(_15986_),
    .ZN(_19298_));
 INV_X1 _37690_ (.A(_15990_),
    .ZN(_16000_));
 INV_X1 _37691_ (.A(_15995_),
    .ZN(_16038_));
 INV_X1 _37692_ (.A(_15999_),
    .ZN(_16039_));
 INV_X1 _37693_ (.A(_16008_),
    .ZN(_16009_));
 INV_X1 _37694_ (.A(_16017_),
    .ZN(_16033_));
 INV_X1 _37695_ (.A(_16024_),
    .ZN(_16065_));
 INV_X1 _37696_ (.A(_16032_),
    .ZN(_16066_));
 INV_X1 _37697_ (.A(_16051_),
    .ZN(_16092_));
 INV_X1 _37698_ (.A(_16056_),
    .ZN(_16093_));
 INV_X1 _37699_ (.A(_16060_),
    .ZN(_16094_));
 INV_X1 _37700_ (.A(_16075_),
    .ZN(_16102_));
 INV_X1 _37701_ (.A(_16079_),
    .ZN(_16117_));
 INV_X1 _37702_ (.A(_16084_),
    .ZN(_16118_));
 INV_X1 _37703_ (.A(_16108_),
    .ZN(_16142_));
 INV_X1 _37704_ (.A(_16112_),
    .ZN(_16143_));
 INV_X1 _37705_ (.A(_16128_),
    .ZN(_16163_));
 INV_X1 _37706_ (.A(_16137_),
    .ZN(_16164_));
 INV_X1 _37707_ (.A(_16149_),
    .ZN(_16158_));
 INV_X1 _37708_ (.A(_16153_),
    .ZN(_16181_));
 INV_X1 _37709_ (.A(_16157_),
    .ZN(_16179_));
 INV_X1 _37710_ (.A(_16187_),
    .ZN(_16188_));
 INV_X1 _37711_ (.A(_16196_),
    .ZN(_19138_));
 INV_X1 _37712_ (.A(_16205_),
    .ZN(_19135_));
 INV_X1 _37713_ (.A(_16213_),
    .ZN(_16215_));
 INV_X1 _37714_ (.A(_16233_),
    .ZN(_16235_));
 INV_X1 _37715_ (.A(_16251_),
    .ZN(_19269_));
 INV_X1 _37716_ (.A(_16260_),
    .ZN(_19273_));
 INV_X1 _37717_ (.A(_16265_),
    .ZN(_16267_));
 INV_X1 _37718_ (.A(_16274_),
    .ZN(_16282_));
 INV_X1 _37719_ (.A(_16279_),
    .ZN(_16281_));
 INV_X1 _37720_ (.A(_16303_),
    .ZN(_16310_));
 INV_X1 _37721_ (.A(_16308_),
    .ZN(_16309_));
 INV_X1 _37722_ (.A(_16324_),
    .ZN(_16338_));
 INV_X1 _37723_ (.A(_16332_),
    .ZN(_16339_));
 INV_X1 _37724_ (.A(_16336_),
    .ZN(_16337_));
 INV_X1 _37725_ (.A(_16352_),
    .ZN(_16366_));
 INV_X1 _37726_ (.A(_16356_),
    .ZN(_16359_));
 INV_X1 _37727_ (.A(_16380_),
    .ZN(_16392_));
 INV_X1 _37728_ (.A(_16387_),
    .ZN(_16393_));
 INV_X1 _37729_ (.A(_16391_),
    .ZN(_16394_));
 INV_X1 _37730_ (.A(_16416_),
    .ZN(_16422_));
 INV_X1 _37731_ (.A(_16421_),
    .ZN(_16423_));
 INV_X1 _37732_ (.A(_16427_),
    .ZN(_16428_));
 INV_X1 _37733_ (.A(_16435_),
    .ZN(_16441_));
 INV_X1 _37734_ (.A(_16439_),
    .ZN(_16440_));
 INV_X1 _37735_ (.A(_16447_),
    .ZN(_16448_));
 INV_X1 _37736_ (.A(_16455_),
    .ZN(_16457_));
 INV_X1 _37737_ (.A(_16468_),
    .ZN(_16470_));
 INV_X1 _37738_ (.A(_16480_),
    .ZN(_16482_));
 INV_X1 _37739_ (.A(_16489_),
    .ZN(_19249_));
 INV_X1 _37740_ (.A(_16492_),
    .ZN(_19248_));
 INV_X1 _37741_ (.A(_16498_),
    .ZN(_19117_));
 INV_X1 _37742_ (.A(_16502_),
    .ZN(_19113_));
 INV_X1 _37743_ (.A(_16506_),
    .ZN(_19114_));
 INV_X1 _37744_ (.A(_16509_),
    .ZN(_16511_));
 INV_X1 _37745_ (.A(_16522_),
    .ZN(_16525_));
 INV_X1 _37746_ (.A(_16532_),
    .ZN(_16534_));
 INV_X1 _37747_ (.A(_16546_),
    .ZN(_19180_));
 INV_X1 _37748_ (.A(_16554_),
    .ZN(_16555_));
 INV_X1 _37749_ (.A(_16567_),
    .ZN(_18708_));
 INV_X1 _37750_ (.A(_16580_),
    .ZN(_16629_));
 INV_X1 _37751_ (.A(_16585_),
    .ZN(_18613_));
 INV_X1 _37752_ (.A(_16588_),
    .ZN(_18614_));
 INV_X1 _37753_ (.A(_16592_),
    .ZN(_18615_));
 INV_X1 _37754_ (.A(_16600_),
    .ZN(_16610_));
 INV_X1 _37755_ (.A(_16609_),
    .ZN(_16611_));
 INV_X1 _37756_ (.A(_16621_),
    .ZN(_17937_));
 INV_X1 _37757_ (.A(_16626_),
    .ZN(_17947_));
 INV_X1 _37758_ (.A(_16638_),
    .ZN(_16648_));
 INV_X1 _37759_ (.A(_16642_),
    .ZN(_18602_));
 INV_X1 _37760_ (.A(_16646_),
    .ZN(_18603_));
 INV_X1 _37761_ (.A(_16661_),
    .ZN(_16667_));
 INV_X1 _37762_ (.A(_16666_),
    .ZN(_16668_));
 INV_X1 _37763_ (.A(_16684_),
    .ZN(_16686_));
 INV_X1 _37764_ (.A(_16701_),
    .ZN(_16710_));
 INV_X1 _37765_ (.A(_16705_),
    .ZN(_16735_));
 INV_X1 _37766_ (.A(_16709_),
    .ZN(_16733_));
 INV_X1 _37767_ (.A(_16726_),
    .ZN(_19160_));
 INV_X1 _37768_ (.A(_16729_),
    .ZN(_19161_));
 INV_X1 _37769_ (.A(_16740_),
    .ZN(_18936_));
 INV_X1 _37770_ (.A(_16744_),
    .ZN(_18937_));
 INV_X1 _37771_ (.A(_16748_),
    .ZN(_18477_));
 INV_X1 _37772_ (.A(_16752_),
    .ZN(_18150_));
 INV_X1 _37773_ (.A(_16768_),
    .ZN(_18467_));
 INV_X1 _37774_ (.A(_16773_),
    .ZN(_18468_));
 INV_X1 _37775_ (.A(_16777_),
    .ZN(_18469_));
 INV_X1 _37776_ (.A(_16785_),
    .ZN(_16795_));
 INV_X1 _37777_ (.A(_16794_),
    .ZN(_16796_));
 INV_X1 _37778_ (.A(_16806_),
    .ZN(_17513_));
 INV_X1 _37779_ (.A(_16811_),
    .ZN(_17530_));
 INV_X1 _37780_ (.A(_16815_),
    .ZN(_17531_));
 INV_X1 _37781_ (.A(_16828_),
    .ZN(_18445_));
 INV_X1 _37782_ (.A(_16837_),
    .ZN(_16844_));
 INV_X1 _37783_ (.A(_16842_),
    .ZN(_16845_));
 INV_X1 _37784_ (.A(_16852_),
    .ZN(_18441_));
 INV_X1 _37785_ (.A(_16856_),
    .ZN(_16866_));
 INV_X1 _37786_ (.A(_16861_),
    .ZN(_18406_));
 INV_X1 _37787_ (.A(_16865_),
    .ZN(_18407_));
 INV_X1 _37788_ (.A(_16874_),
    .ZN(_16875_));
 INV_X1 _37789_ (.A(_16883_),
    .ZN(_18409_));
 INV_X1 _37790_ (.A(_16894_),
    .ZN(_18102_));
 INV_X1 _37791_ (.A(_16898_),
    .ZN(_18103_));
 INV_X1 _37792_ (.A(_16912_),
    .ZN(_18387_));
 INV_X1 _37793_ (.A(_16917_),
    .ZN(_18388_));
 INV_X1 _37794_ (.A(_16926_),
    .ZN(_16939_));
 INV_X1 _37795_ (.A(_16934_),
    .ZN(_16940_));
 INV_X1 _37796_ (.A(_16938_),
    .ZN(_16941_));
 INV_X1 _37797_ (.A(_16948_),
    .ZN(_18384_));
 INV_X1 _37798_ (.A(_16952_),
    .ZN(_17567_));
 INV_X1 _37799_ (.A(_16956_),
    .ZN(_17568_));
 INV_X1 _37800_ (.A(_16965_),
    .ZN(_18911_));
 INV_X1 _37801_ (.A(_16974_),
    .ZN(_18371_));
 INV_X1 _37802_ (.A(_16979_),
    .ZN(_18844_));
 INV_X1 _37803_ (.A(_16983_),
    .ZN(_18845_));
 INV_X1 _37804_ (.A(_16987_),
    .ZN(_18578_));
 INV_X1 _37805_ (.A(_16991_),
    .ZN(_18049_));
 INV_X1 _37806_ (.A(_17007_),
    .ZN(_18565_));
 INV_X1 _37807_ (.A(_17012_),
    .ZN(_18566_));
 INV_X1 _37808_ (.A(_17016_),
    .ZN(_18567_));
 INV_X1 _37809_ (.A(_17024_),
    .ZN(_17034_));
 INV_X1 _37810_ (.A(_17033_),
    .ZN(_17035_));
 INV_X1 _37811_ (.A(_17049_),
    .ZN(_17577_));
 INV_X1 _37812_ (.A(_17054_),
    .ZN(_17576_));
 INV_X1 _37813_ (.A(_17062_),
    .ZN(_17073_));
 INV_X1 _37814_ (.A(_17072_),
    .ZN(_17074_));
 INV_X1 _37815_ (.A(_17081_),
    .ZN(_17090_));
 INV_X1 _37816_ (.A(_17085_),
    .ZN(_18548_));
 INV_X1 _37817_ (.A(_17089_),
    .ZN(_18550_));
 INV_X1 _37818_ (.A(_17108_),
    .ZN(_17109_));
 INV_X1 _37819_ (.A(_17117_),
    .ZN(_18795_));
 INV_X1 _37820_ (.A(_17121_),
    .ZN(_18796_));
 INV_X1 _37821_ (.A(_17124_),
    .ZN(_18526_));
 INV_X1 _37822_ (.A(_17128_),
    .ZN(_17624_));
 INV_X1 _37823_ (.A(_17136_),
    .ZN(_17142_));
 INV_X1 _37824_ (.A(_17141_),
    .ZN(_17143_));
 INV_X1 _37825_ (.A(_17158_),
    .ZN(_17190_));
 INV_X1 _37826_ (.A(_17163_),
    .ZN(_18514_));
 INV_X1 _37827_ (.A(_17166_),
    .ZN(_18513_));
 INV_X1 _37828_ (.A(_17170_),
    .ZN(_18515_));
 INV_X1 _37829_ (.A(_17187_),
    .ZN(_18000_));
 INV_X1 _37830_ (.A(_17199_),
    .ZN(_17210_));
 INV_X1 _37831_ (.A(_17209_),
    .ZN(_17211_));
 INV_X1 _37832_ (.A(_17223_),
    .ZN(_18500_));
 INV_X1 _37833_ (.A(_17228_),
    .ZN(_18501_));
 INV_X1 _37834_ (.A(_17246_),
    .ZN(_17248_));
 INV_X1 _37835_ (.A(_17256_),
    .ZN(_17265_));
 INV_X1 _37836_ (.A(_17260_),
    .ZN(_18657_));
 INV_X1 _37837_ (.A(_17264_),
    .ZN(_18659_));
 INV_X1 _37838_ (.A(_17274_),
    .ZN(_17285_));
 INV_X1 _37839_ (.A(_17284_),
    .ZN(_17286_));
 INV_X1 _37840_ (.A(_17301_),
    .ZN(_17309_));
 INV_X1 _37841_ (.A(_17315_),
    .ZN(_18665_));
 INV_X1 _37842_ (.A(_17319_),
    .ZN(_18664_));
 INV_X1 _37843_ (.A(_17331_),
    .ZN(_17341_));
 INV_X1 _37844_ (.A(_17336_),
    .ZN(_17342_));
 INV_X1 _37845_ (.A(_17352_),
    .ZN(_18751_));
 INV_X1 _37846_ (.A(_17356_),
    .ZN(_18752_));
 INV_X1 _37847_ (.A(_17360_),
    .ZN(_18682_));
 INV_X1 _37848_ (.A(_17364_),
    .ZN(_17385_));
 INV_X1 _37849_ (.A(_17369_),
    .ZN(_17371_));
 INV_X1 _37850_ (.A(_17378_),
    .ZN(_18773_));
 INV_X1 _37851_ (.A(_17392_),
    .ZN(_17402_));
 INV_X1 _37852_ (.A(_17397_),
    .ZN(_18673_));
 INV_X1 _37853_ (.A(_17401_),
    .ZN(_18674_));
 INV_X1 _37854_ (.A(_17410_),
    .ZN(_18676_));
 INV_X1 _37855_ (.A(_17417_),
    .ZN(_17974_));
 INV_X1 _37856_ (.A(_17425_),
    .ZN(_17975_));
 INV_X1 _37857_ (.A(_17435_),
    .ZN(_17437_));
 INV_X1 _37858_ (.A(_17453_),
    .ZN(_17502_));
 INV_X1 _37859_ (.A(_17458_),
    .ZN(_18298_));
 INV_X1 _37860_ (.A(_17462_),
    .ZN(_18299_));
 INV_X1 _37861_ (.A(_17474_),
    .ZN(_17486_));
 INV_X1 _37862_ (.A(_17481_),
    .ZN(_17487_));
 INV_X1 _37863_ (.A(_17485_),
    .ZN(_17488_));
 INV_X1 _37864_ (.A(_17499_),
    .ZN(_17885_));
 INV_X1 _37865_ (.A(_17507_),
    .ZN(_17884_));
 INV_X1 _37866_ (.A(_17521_),
    .ZN(_18462_));
 INV_X1 _37867_ (.A(_17525_),
    .ZN(_18463_));
 INV_X1 _37868_ (.A(_17542_),
    .ZN(_18455_));
 INV_X1 _37869_ (.A(_17551_),
    .ZN(_18456_));
 INV_X1 _37870_ (.A(_17575_),
    .ZN(_18377_));
 INV_X1 _37871_ (.A(_17588_),
    .ZN(_18557_));
 INV_X1 _37872_ (.A(_17593_),
    .ZN(_18556_));
 INV_X1 _37873_ (.A(_17597_),
    .ZN(_18558_));
 INV_X1 _37874_ (.A(_17608_),
    .ZN(_17618_));
 INV_X1 _37875_ (.A(_17613_),
    .ZN(_18522_));
 INV_X1 _37876_ (.A(_17617_),
    .ZN(_18523_));
 INV_X1 _37877_ (.A(_17629_),
    .ZN(_18519_));
 INV_X1 _37878_ (.A(_17634_),
    .ZN(_17636_));
 INV_X1 _37879_ (.A(_17643_),
    .ZN(_17649_));
 INV_X1 _37880_ (.A(_17647_),
    .ZN(_18630_));
 INV_X1 _37881_ (.A(_17660_),
    .ZN(_18626_));
 INV_X1 _37882_ (.A(_17665_),
    .ZN(_18622_));
 INV_X1 _37883_ (.A(_17669_),
    .ZN(_18623_));
 INV_X1 _37884_ (.A(_17674_),
    .ZN(_19025_));
 INV_X1 _37885_ (.A(_17678_),
    .ZN(_19024_));
 INV_X1 _37886_ (.A(_17682_),
    .ZN(_18364_));
 INV_X1 _37887_ (.A(_17686_),
    .ZN(_18253_));
 INV_X1 _37888_ (.A(_17690_),
    .ZN(_17700_));
 INV_X1 _37889_ (.A(_17699_),
    .ZN(_17701_));
 INV_X1 _37890_ (.A(_17719_),
    .ZN(_18351_));
 INV_X1 _37891_ (.A(_17724_),
    .ZN(_18350_));
 INV_X1 _37892_ (.A(_17728_),
    .ZN(_18349_));
 INV_X1 _37893_ (.A(_17744_),
    .ZN(_17753_));
 INV_X1 _37894_ (.A(_17749_),
    .ZN(_17754_));
 INV_X1 _37895_ (.A(_17765_),
    .ZN(_18342_));
 INV_X1 _37896_ (.A(_17770_),
    .ZN(_18343_));
 INV_X1 _37897_ (.A(_17774_),
    .ZN(_18344_));
 INV_X1 _37898_ (.A(_17787_),
    .ZN(_18196_));
 INV_X1 _37899_ (.A(_17796_),
    .ZN(_18197_));
 INV_X1 _37900_ (.A(_17805_),
    .ZN(_19046_));
 INV_X1 _37901_ (.A(_17810_),
    .ZN(_17812_));
 INV_X1 _37902_ (.A(_17828_),
    .ZN(_17835_));
 INV_X1 _37903_ (.A(_17832_),
    .ZN(_17833_));
 INV_X1 _37904_ (.A(_17841_),
    .ZN(_17852_));
 INV_X1 _37905_ (.A(_17847_),
    .ZN(_18303_));
 INV_X1 _37906_ (.A(_17851_),
    .ZN(_18304_));
 INV_X1 _37907_ (.A(_17874_),
    .ZN(_18294_));
 INV_X1 _37908_ (.A(_17879_),
    .ZN(_18293_));
 INV_X1 _37909_ (.A(_17892_),
    .ZN(_18290_));
 INV_X1 _37910_ (.A(_17896_),
    .ZN(_17917_));
 INV_X1 _37911_ (.A(_17900_),
    .ZN(_17915_));
 INV_X1 _37912_ (.A(_17910_),
    .ZN(_18288_));
 INV_X1 _37913_ (.A(_17924_),
    .ZN(_18283_));
 INV_X1 _37914_ (.A(_17934_),
    .ZN(_18609_));
 INV_X1 _37915_ (.A(_17942_),
    .ZN(_18608_));
 INV_X1 _37916_ (.A(_17960_),
    .ZN(_18669_));
 INV_X1 _37917_ (.A(_17965_),
    .ZN(_18670_));
 INV_X1 _37918_ (.A(_17969_),
    .ZN(_18671_));
 INV_X1 _37919_ (.A(_17984_),
    .ZN(_18822_));
 INV_X1 _37920_ (.A(_17989_),
    .ZN(_17991_));
 INV_X1 _37921_ (.A(_18012_),
    .ZN(_18508_));
 INV_X1 _37922_ (.A(_18016_),
    .ZN(_18507_));
 INV_X1 _37923_ (.A(_18020_),
    .ZN(_18509_));
 INV_X1 _37924_ (.A(_18031_),
    .ZN(_18867_));
 INV_X1 _37925_ (.A(_18036_),
    .ZN(_18037_));
 INV_X1 _37926_ (.A(_18055_),
    .ZN(_18065_));
 INV_X1 _37927_ (.A(_18060_),
    .ZN(_18569_));
 INV_X1 _37928_ (.A(_18064_),
    .ZN(_18570_));
 INV_X1 _37929_ (.A(_18071_),
    .ZN(_18572_));
 INV_X1 _37930_ (.A(_18080_),
    .ZN(_18117_));
 INV_X1 _37931_ (.A(_18090_),
    .ZN(_18403_));
 INV_X1 _37932_ (.A(_18093_),
    .ZN(_18402_));
 INV_X1 _37933_ (.A(_18097_),
    .ZN(_18404_));
 INV_X1 _37934_ (.A(_18114_),
    .ZN(_18397_));
 INV_X1 _37935_ (.A(_18126_),
    .ZN(_18129_));
 INV_X1 _37936_ (.A(_18135_),
    .ZN(_18145_));
 INV_X1 _37937_ (.A(_18140_),
    .ZN(_18474_));
 INV_X1 _37938_ (.A(_18144_),
    .ZN(_18475_));
 INV_X1 _37939_ (.A(_18156_),
    .ZN(_18471_));
 INV_X1 _37940_ (.A(_18165_),
    .ZN(_19000_));
 INV_X1 _37941_ (.A(_18174_),
    .ZN(_18278_));
 INV_X1 _37942_ (.A(_18182_),
    .ZN(_18188_));
 INV_X1 _37943_ (.A(_18186_),
    .ZN(_18307_));
 INV_X1 _37944_ (.A(_18195_),
    .ZN(_18311_));
 INV_X1 _37945_ (.A(_18204_),
    .ZN(_18214_));
 INV_X1 _37946_ (.A(_18208_),
    .ZN(_18334_));
 INV_X1 _37947_ (.A(_18212_),
    .ZN(_18336_));
 INV_X1 _37948_ (.A(_18226_),
    .ZN(_18228_));
 INV_X1 _37949_ (.A(_18235_),
    .ZN(_18729_));
 INV_X1 _37950_ (.A(_18244_),
    .ZN(_18890_));
 INV_X1 _37951_ (.A(_18248_),
    .ZN(_18889_));
 INV_X1 _37952_ (.A(_18251_),
    .ZN(_18413_));
 INV_X1 _37953_ (.A(_18260_),
    .ZN(_18270_));
 INV_X1 _37954_ (.A(_18265_),
    .ZN(_18355_));
 INV_X1 _37955_ (.A(_18269_),
    .ZN(_18356_));
 INV_X1 _37956_ (.A(_18276_),
    .ZN(_18358_));
 INV_X1 _37957_ (.A(_18318_),
    .ZN(_18982_));
 INV_X1 _37958_ (.A(_18321_),
    .ZN(_18983_));
 INV_X1 _37959_ (.A(_18333_),
    .ZN(_19042_));
 INV_X1 _37960_ (.A(_18383_),
    .ZN(_18914_));
 INV_X1 _37961_ (.A(_18422_),
    .ZN(_18893_));
 INV_X1 _37962_ (.A(_18435_),
    .ZN(_18958_));
 INV_X1 _37963_ (.A(_18451_),
    .ZN(_18452_));
 INV_X1 _37964_ (.A(_18486_),
    .ZN(_18940_));
 INV_X1 _37965_ (.A(_18498_),
    .ZN(_18819_));
 INV_X1 _37966_ (.A(_18535_),
    .ZN(_18800_));
 INV_X1 _37967_ (.A(_18547_),
    .ZN(_18864_));
 INV_X1 _37968_ (.A(_18592_),
    .ZN(_18726_));
 INV_X1 _37969_ (.A(_18618_),
    .ZN(_18619_));
 INV_X1 _37970_ (.A(_18636_),
    .ZN(_18703_));
 INV_X1 _37971_ (.A(_18640_),
    .ZN(_18704_));
 INV_X1 _37972_ (.A(_18648_),
    .ZN(_18770_));
 INV_X1 _37973_ (.A(_18690_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[10] ));
 INV_X1 _37974_ (.A(_18692_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[11] ));
 INV_X1 _37975_ (.A(_18694_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[12] ));
 INV_X1 _37976_ (.A(_18696_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[13] ));
 INV_X1 _37977_ (.A(_18698_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[14] ));
 INV_X1 _37978_ (.A(_18700_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[15] ));
 INV_X1 _37979_ (.A(_18702_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[16] ));
 INV_X1 _37980_ (.A(_18706_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[17] ));
 INV_X1 _37981_ (.A(_18711_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[18] ));
 INV_X1 _37982_ (.A(_18716_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[19] ));
 INV_X1 _37983_ (.A(_18725_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[5] ));
 INV_X1 _37984_ (.A(_18728_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[6] ));
 INV_X1 _37985_ (.A(_18732_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[7] ));
 INV_X1 _37986_ (.A(_18734_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[8] ));
 INV_X1 _37987_ (.A(_18736_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[9] ));
 INV_X1 _37988_ (.A(_18738_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[10] ));
 INV_X1 _37989_ (.A(_18740_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[11] ));
 INV_X1 _37990_ (.A(_18742_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[12] ));
 INV_X1 _37991_ (.A(_18744_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[13] ));
 INV_X1 _37992_ (.A(_18746_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[14] ));
 INV_X1 _37993_ (.A(_18748_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[15] ));
 INV_X1 _37994_ (.A(_18750_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[16] ));
 INV_X1 _37995_ (.A(_18754_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[17] ));
 INV_X1 _37996_ (.A(_18760_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[19] ));
 INV_X1 _37997_ (.A(_18769_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[5] ));
 INV_X1 _37998_ (.A(_18772_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[6] ));
 INV_X1 _37999_ (.A(_18776_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[7] ));
 INV_X1 _38000_ (.A(_18778_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[8] ));
 INV_X1 _38001_ (.A(_18780_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[9] ));
 INV_X1 _38002_ (.A(_18782_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[10] ));
 INV_X1 _38003_ (.A(_18784_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[11] ));
 INV_X1 _38004_ (.A(_18786_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[12] ));
 INV_X1 _38005_ (.A(_18788_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[13] ));
 INV_X1 _38006_ (.A(_18790_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[14] ));
 INV_X1 _38007_ (.A(_18792_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[15] ));
 INV_X1 _38008_ (.A(_18794_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[16] ));
 INV_X1 _38009_ (.A(_18798_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[17] ));
 INV_X1 _38010_ (.A(_18803_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[18] ));
 INV_X1 _38011_ (.A(_18808_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[19] ));
 INV_X1 _38012_ (.A(_18817_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[5] ));
 INV_X1 _38013_ (.A(_18821_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[6] ));
 INV_X1 _38014_ (.A(_18825_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[7] ));
 INV_X1 _38015_ (.A(_18827_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[8] ));
 INV_X1 _38016_ (.A(_18829_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[9] ));
 INV_X1 _38017_ (.A(_18831_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[10] ));
 INV_X1 _38018_ (.A(_18833_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[11] ));
 INV_X1 _38019_ (.A(_18835_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[12] ));
 INV_X1 _38020_ (.A(_18837_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[13] ));
 INV_X1 _38021_ (.A(_18839_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[14] ));
 INV_X1 _38022_ (.A(_18841_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[15] ));
 INV_X1 _38023_ (.A(_18843_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[16] ));
 INV_X1 _38024_ (.A(_18847_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[17] ));
 INV_X1 _38025_ (.A(_18853_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[19] ));
 INV_X1 _38026_ (.A(_18862_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[5] ));
 INV_X1 _38027_ (.A(_18866_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[6] ));
 INV_X1 _38028_ (.A(_18870_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[7] ));
 INV_X1 _38029_ (.A(_18872_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[8] ));
 INV_X1 _38030_ (.A(_18874_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[9] ));
 INV_X1 _38031_ (.A(_18876_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[10] ));
 INV_X1 _38032_ (.A(_18878_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[11] ));
 INV_X1 _38033_ (.A(_18880_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[12] ));
 INV_X1 _38034_ (.A(_18882_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[13] ));
 INV_X1 _38035_ (.A(_18884_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[14] ));
 INV_X1 _38036_ (.A(_18886_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[15] ));
 INV_X1 _38037_ (.A(_18888_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[16] ));
 INV_X1 _38038_ (.A(_18892_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[17] ));
 INV_X1 _38039_ (.A(_18897_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[18] ));
 INV_X1 _38040_ (.A(_18901_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[19] ));
 INV_X1 _38041_ (.A(_18910_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[5] ));
 INV_X1 _38042_ (.A(_18913_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[6] ));
 INV_X1 _38043_ (.A(_18917_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[7] ));
 INV_X1 _38044_ (.A(_18919_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[8] ));
 INV_X1 _38045_ (.A(_18921_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[9] ));
 INV_X1 _38046_ (.A(_18923_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[10] ));
 INV_X1 _38047_ (.A(_18925_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[11] ));
 INV_X1 _38048_ (.A(_18927_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[12] ));
 INV_X1 _38049_ (.A(_18929_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[13] ));
 INV_X1 _38050_ (.A(_18931_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[14] ));
 INV_X1 _38051_ (.A(_18933_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[15] ));
 INV_X1 _38052_ (.A(_18935_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[16] ));
 INV_X1 _38053_ (.A(_18939_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[17] ));
 INV_X1 _38054_ (.A(_18944_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[18] ));
 INV_X1 _38055_ (.A(_18948_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[19] ));
 INV_X1 _38056_ (.A(_18957_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[5] ));
 INV_X1 _38057_ (.A(_18960_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[6] ));
 INV_X1 _38058_ (.A(_18963_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[7] ));
 INV_X1 _38059_ (.A(_18965_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[8] ));
 INV_X1 _38060_ (.A(_18967_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[9] ));
 INV_X1 _38061_ (.A(_18969_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[10] ));
 INV_X1 _38062_ (.A(_18971_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[11] ));
 INV_X1 _38063_ (.A(_18973_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[12] ));
 INV_X1 _38064_ (.A(_18975_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[13] ));
 INV_X1 _38065_ (.A(_18977_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[14] ));
 INV_X1 _38066_ (.A(_18979_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[15] ));
 INV_X1 _38067_ (.A(_18981_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[16] ));
 INV_X1 _38068_ (.A(_18985_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[17] ));
 INV_X1 _38069_ (.A(_18990_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[19] ));
 INV_X1 _38070_ (.A(_18999_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[5] ));
 INV_X1 _38071_ (.A(_19002_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[6] ));
 INV_X1 _38072_ (.A(_19005_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[7] ));
 INV_X1 _38073_ (.A(_19007_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[8] ));
 INV_X1 _38074_ (.A(_19009_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[9] ));
 INV_X1 _38075_ (.A(_19011_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[10] ));
 INV_X1 _38076_ (.A(_19013_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[11] ));
 INV_X1 _38077_ (.A(_19015_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[12] ));
 INV_X1 _38078_ (.A(_19017_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[13] ));
 INV_X1 _38079_ (.A(_19019_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[14] ));
 INV_X1 _38080_ (.A(_19021_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[15] ));
 INV_X1 _38081_ (.A(_19023_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[16] ));
 INV_X1 _38082_ (.A(_19027_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[17] ));
 INV_X1 _38083_ (.A(_19032_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[19] ));
 INV_X1 _38084_ (.A(_19041_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[5] ));
 INV_X1 _38085_ (.A(_19044_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[6] ));
 INV_X1 _38086_ (.A(_19048_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[7] ));
 INV_X1 _38087_ (.A(_19050_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[8] ));
 INV_X1 _38088_ (.A(_19052_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[9] ));
 INV_X1 _38089_ (.A(_19054_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[10] ));
 INV_X1 _38090_ (.A(_19056_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[11] ));
 INV_X1 _38091_ (.A(_19058_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[12] ));
 INV_X1 _38092_ (.A(_19060_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[13] ));
 INV_X1 _38093_ (.A(_19062_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[14] ));
 INV_X1 _38094_ (.A(_19064_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[15] ));
 INV_X1 _38095_ (.A(_19066_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[16] ));
 INV_X1 _38096_ (.A(_19070_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[17] ));
 INV_X1 _38097_ (.A(_19075_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[19] ));
 INV_X1 _38098_ (.A(_19080_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[3] ));
 INV_X1 _38099_ (.A(_19086_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[5] ));
 INV_X1 _38100_ (.A(_19090_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[6] ));
 INV_X1 _38101_ (.A(_19094_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[7] ));
 INV_X1 _38102_ (.A(_19096_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[8] ));
 INV_X1 _38103_ (.A(_19098_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[9] ));
 INV_X1 _38104_ (.A(_19100_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[10] ));
 INV_X1 _38105_ (.A(_19102_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[11] ));
 INV_X1 _38106_ (.A(_19104_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[12] ));
 INV_X1 _38107_ (.A(_19106_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[13] ));
 INV_X1 _38108_ (.A(_19108_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[14] ));
 INV_X1 _38109_ (.A(_19110_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[15] ));
 INV_X1 _38110_ (.A(_19112_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[16] ));
 INV_X1 _38111_ (.A(_19116_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[17] ));
 INV_X1 _38112_ (.A(_19121_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[18] ));
 INV_X1 _38113_ (.A(_19125_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[19] ));
 INV_X1 _38114_ (.A(_19134_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[5] ));
 INV_X1 _38115_ (.A(_19137_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[6] ));
 INV_X1 _38116_ (.A(_19141_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[7] ));
 INV_X1 _38117_ (.A(_19143_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[8] ));
 INV_X1 _38118_ (.A(_19145_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[9] ));
 INV_X1 _38119_ (.A(_19147_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[10] ));
 INV_X1 _38120_ (.A(_19149_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[11] ));
 INV_X1 _38121_ (.A(_19151_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[12] ));
 INV_X1 _38122_ (.A(_19153_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[13] ));
 INV_X1 _38123_ (.A(_19155_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[14] ));
 INV_X1 _38124_ (.A(_19157_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[15] ));
 INV_X1 _38125_ (.A(_19159_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[16] ));
 INV_X1 _38126_ (.A(_19163_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[17] ));
 INV_X1 _38127_ (.A(_19168_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[19] ));
 INV_X1 _38128_ (.A(_19173_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[3] ));
 INV_X1 _38129_ (.A(_19179_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[5] ));
 INV_X1 _38130_ (.A(_19182_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[6] ));
 INV_X1 _38131_ (.A(_19185_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[7] ));
 INV_X1 _38132_ (.A(_19187_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[8] ));
 INV_X1 _38133_ (.A(_19189_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[9] ));
 INV_X1 _38134_ (.A(_19191_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[10] ));
 INV_X1 _38135_ (.A(_19193_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[11] ));
 INV_X1 _38136_ (.A(_19195_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[12] ));
 INV_X1 _38137_ (.A(_19197_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[13] ));
 INV_X1 _38138_ (.A(_19199_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[14] ));
 INV_X1 _38139_ (.A(_19201_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[15] ));
 INV_X1 _38140_ (.A(_19203_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[16] ));
 INV_X1 _38141_ (.A(_19207_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[17] ));
 INV_X1 _38142_ (.A(_19212_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[19] ));
 INV_X1 _38143_ (.A(_19217_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[3] ));
 INV_X1 _38144_ (.A(_19223_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[5] ));
 INV_X1 _38145_ (.A(_19226_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[6] ));
 INV_X1 _38146_ (.A(_19229_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[7] ));
 INV_X1 _38147_ (.A(_19231_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[8] ));
 INV_X1 _38148_ (.A(_19233_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[9] ));
 INV_X1 _38149_ (.A(_19235_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[10] ));
 INV_X1 _38150_ (.A(_19237_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[11] ));
 INV_X1 _38151_ (.A(_19239_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[12] ));
 INV_X1 _38152_ (.A(_19241_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[13] ));
 INV_X1 _38153_ (.A(_19243_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[14] ));
 INV_X1 _38154_ (.A(_19245_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[15] ));
 INV_X1 _38155_ (.A(_19247_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[16] ));
 INV_X1 _38156_ (.A(_19251_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[17] ));
 INV_X1 _38157_ (.A(_19256_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[19] ));
 INV_X1 _38158_ (.A(_19261_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[3] ));
 INV_X1 _38159_ (.A(_19267_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[5] ));
 INV_X1 _38160_ (.A(_19271_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[6] ));
 INV_X1 _38161_ (.A(_19275_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[7] ));
 INV_X1 _38162_ (.A(_19277_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[8] ));
 INV_X1 _38163_ (.A(_19279_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[9] ));
 INV_X1 _38164_ (.A(_19281_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[10] ));
 INV_X1 _38165_ (.A(_19283_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[11] ));
 INV_X1 _38166_ (.A(_19285_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[12] ));
 INV_X1 _38167_ (.A(_19287_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[13] ));
 INV_X1 _38168_ (.A(_19289_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[14] ));
 INV_X1 _38169_ (.A(_19291_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[15] ));
 INV_X1 _38170_ (.A(_19293_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[16] ));
 INV_X1 _38171_ (.A(_19297_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[17] ));
 INV_X1 _38172_ (.A(_19302_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[18] ));
 INV_X1 _38173_ (.A(_19306_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[19] ));
 INV_X1 _38174_ (.A(_19311_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[3] ));
 INV_X1 _38175_ (.A(_19317_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[5] ));
 INV_X1 _38176_ (.A(_19321_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[6] ));
 INV_X1 _38177_ (.A(_19325_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[7] ));
 INV_X1 _38178_ (.A(_19327_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[8] ));
 INV_X1 _38179_ (.A(_19329_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[9] ));
 INV_X1 _38180_ (.A(_19331_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[10] ));
 INV_X1 _38181_ (.A(_19333_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[11] ));
 INV_X1 _38182_ (.A(_19335_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[12] ));
 INV_X1 _38183_ (.A(_19337_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[13] ));
 INV_X1 _38184_ (.A(_19339_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[14] ));
 INV_X1 _38185_ (.A(_19341_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[15] ));
 INV_X1 _38186_ (.A(_19343_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[16] ));
 INV_X1 _38187_ (.A(_19347_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[17] ));
 INV_X1 _38188_ (.A(_19352_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[18] ));
 INV_X1 _38189_ (.A(_19356_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[19] ));
 INV_X1 _38190_ (.A(_19361_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[3] ));
 INV_X1 _38191_ (.A(_19367_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[5] ));
 INV_X1 _38192_ (.A(_19370_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[6] ));
 INV_X1 _38193_ (.A(_19373_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[7] ));
 INV_X1 _38194_ (.A(_19375_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[8] ));
 INV_X1 _38195_ (.A(_19377_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[9] ));
 INV_X1 _38196_ (.A(_19379_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[10] ));
 INV_X1 _38197_ (.A(_19381_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[11] ));
 INV_X1 _38198_ (.A(_19383_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[12] ));
 INV_X1 _38199_ (.A(_19385_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[13] ));
 INV_X1 _38200_ (.A(_19387_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[14] ));
 INV_X1 _38201_ (.A(_19389_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[15] ));
 INV_X1 _38202_ (.A(_19391_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[16] ));
 INV_X1 _38203_ (.A(_19395_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[17] ));
 INV_X1 _38204_ (.A(_19400_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[19] ));
 INV_X1 _38205_ (.A(_19405_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[3] ));
 INV_X1 _38206_ (.A(_19411_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[5] ));
 INV_X1 _38207_ (.A(_19415_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[6] ));
 INV_X1 _38208_ (.A(_19419_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[7] ));
 INV_X1 _38209_ (.A(_19421_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[8] ));
 INV_X1 _38210_ (.A(_19423_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[9] ));
 INV_X1 _38211_ (.A(_14530_),
    .ZN(_14990_));
 INV_X1 _38212_ (.A(_14535_),
    .ZN(_14991_));
 INV_X1 _38213_ (.A(_14549_),
    .ZN(_14542_));
 INV_X1 _38214_ (.A(_14554_),
    .ZN(_14543_));
 INV_X1 _38215_ (.A(_14567_),
    .ZN(_14562_));
 INV_X1 _38216_ (.A(_14572_),
    .ZN(_19208_));
 INV_X1 _38217_ (.A(_14584_),
    .ZN(_15346_));
 INV_X1 _38218_ (.A(_14597_),
    .ZN(_14590_));
 INV_X1 _38219_ (.A(_14601_),
    .ZN(_14591_));
 INV_X1 _38220_ (.A(_14611_),
    .ZN(_14604_));
 INV_X1 _38221_ (.A(_14614_),
    .ZN(_19210_));
 INV_X1 _38222_ (.A(_14622_),
    .ZN(_19092_));
 INV_X1 _38223_ (.A(_14636_),
    .ZN(_19084_));
 INV_X1 _38224_ (.A(_14640_),
    .ZN(_14678_));
 INV_X1 _38225_ (.A(_14650_),
    .ZN(_14643_));
 INV_X1 _38226_ (.A(_14658_),
    .ZN(_14642_));
 INV_X1 _38227_ (.A(_14667_),
    .ZN(_15128_));
 INV_X1 _38228_ (.A(_14675_),
    .ZN(_15129_));
 INV_X1 _38229_ (.A(_14693_),
    .ZN(_14686_));
 INV_X1 _38230_ (.A(_14702_),
    .ZN(_14688_));
 INV_X1 _38231_ (.A(_14707_),
    .ZN(_19409_));
 INV_X1 _38232_ (.A(_14727_),
    .ZN(_14747_));
 INV_X1 _38233_ (.A(_14730_),
    .ZN(_19417_));
 INV_X1 _38234_ (.A(_14735_),
    .ZN(_14765_));
 INV_X1 _38235_ (.A(_14739_),
    .ZN(_14771_));
 INV_X1 _38236_ (.A(_14744_),
    .ZN(_14770_));
 INV_X1 _38237_ (.A(_14777_),
    .ZN(_14822_));
 INV_X1 _38238_ (.A(_14787_),
    .ZN(_14821_));
 INV_X1 _38239_ (.A(_14794_),
    .ZN(_14825_));
 INV_X1 _38240_ (.A(_14801_),
    .ZN(_14843_));
 INV_X1 _38241_ (.A(_14805_),
    .ZN(_14851_));
 INV_X1 _38242_ (.A(_14810_),
    .ZN(_14850_));
 INV_X1 _38243_ (.A(_14814_),
    .ZN(_14852_));
 INV_X1 _38244_ (.A(_14834_),
    .ZN(_14879_));
 INV_X1 _38245_ (.A(_14839_),
    .ZN(_14878_));
 INV_X1 _38246_ (.A(_14860_),
    .ZN(_14902_));
 INV_X1 _38247_ (.A(_14864_),
    .ZN(_14889_));
 INV_X1 _38248_ (.A(_14867_),
    .ZN(_14903_));
 INV_X1 _38249_ (.A(_14871_),
    .ZN(_14904_));
 INV_X1 _38250_ (.A(_14912_),
    .ZN(_14933_));
 INV_X1 _38251_ (.A(_14916_),
    .ZN(_14931_));
 INV_X1 _38252_ (.A(_14922_),
    .ZN(_14941_));
 INV_X1 _38253_ (.A(_14929_),
    .ZN(_14945_));
 INV_X1 _38254_ (.A(_14938_),
    .ZN(_14954_));
 INV_X1 _38255_ (.A(_14960_),
    .ZN(_19396_));
 INV_X1 _38256_ (.A(_14966_),
    .ZN(_19398_));
 INV_X1 _38257_ (.A(_14971_),
    .ZN(_15338_));
 INV_X1 _38258_ (.A(_14975_),
    .ZN(_15315_));
 INV_X1 _38259_ (.A(_14979_),
    .ZN(_15339_));
 INV_X1 _38260_ (.A(_14983_),
    .ZN(_15340_));
 INV_X1 _38261_ (.A(_14999_),
    .ZN(_15046_));
 INV_X1 _38262_ (.A(_15017_),
    .ZN(_15043_));
 INV_X1 _38263_ (.A(_15027_),
    .ZN(_15042_));
 INV_X1 _38264_ (.A(_15040_),
    .ZN(_15035_));
 INV_X1 _38265_ (.A(_15052_),
    .ZN(_15072_));
 INV_X1 _38266_ (.A(_15056_),
    .ZN(_15090_));
 INV_X1 _38267_ (.A(_15065_),
    .ZN(_15071_));
 INV_X1 _38268_ (.A(_15083_),
    .ZN(_15098_));
 INV_X1 _38269_ (.A(_15088_),
    .ZN(_15099_));
 INV_X1 _38270_ (.A(_15106_),
    .ZN(_15177_));
 INV_X1 _38271_ (.A(_15109_),
    .ZN(_15191_));
 INV_X1 _38272_ (.A(_15114_),
    .ZN(_15189_));
 INV_X1 _38273_ (.A(_15118_),
    .ZN(_15190_));
 INV_X1 _38274_ (.A(_15126_),
    .ZN(_19073_));
 INV_X1 _38275_ (.A(_15137_),
    .ZN(_15406_));
 INV_X1 _38276_ (.A(_15141_),
    .ZN(_15414_));
 INV_X1 _38277_ (.A(_15144_),
    .ZN(_15405_));
 INV_X1 _38278_ (.A(_15148_),
    .ZN(_15407_));
 INV_X1 _38279_ (.A(_15158_),
    .ZN(_19071_));
 INV_X1 _38280_ (.A(_15170_),
    .ZN(_15198_));
 INV_X1 _38281_ (.A(_15207_),
    .ZN(_15201_));
 INV_X1 _38282_ (.A(_15212_),
    .ZN(_15220_));
 INV_X1 _38283_ (.A(_15216_),
    .ZN(_15219_));
 INV_X1 _38284_ (.A(_15229_),
    .ZN(_15240_));
 INV_X1 _38285_ (.A(_15233_),
    .ZN(_15223_));
 INV_X1 _38286_ (.A(_15250_),
    .ZN(_15319_));
 INV_X1 _38287_ (.A(_15254_),
    .ZN(_15318_));
 INV_X1 _38288_ (.A(_15260_),
    .ZN(_15326_));
 INV_X1 _38289_ (.A(_15284_),
    .ZN(_15275_));
 INV_X1 _38290_ (.A(_15287_),
    .ZN(_15273_));
 INV_X1 _38291_ (.A(_15291_),
    .ZN(_15274_));
 INV_X1 _38292_ (.A(_15307_),
    .ZN(_15301_));
 INV_X1 _38293_ (.A(_15324_),
    .ZN(_15349_));
 INV_X1 _38294_ (.A(_15356_),
    .ZN(_19365_));
 INV_X1 _38295_ (.A(_15371_),
    .ZN(_19221_));
 INV_X1 _38296_ (.A(_15376_),
    .ZN(_15391_));
 INV_X1 _38297_ (.A(_15379_),
    .ZN(_19371_));
 INV_X1 _38298_ (.A(_15389_),
    .ZN(_15435_));
 INV_X1 _38299_ (.A(_15398_),
    .ZN(_15432_));
 INV_X1 _38300_ (.A(_15454_),
    .ZN(_15492_));
 INV_X1 _38301_ (.A(_15467_),
    .ZN(_15488_));
 INV_X1 _38302_ (.A(_15472_),
    .ZN(_15489_));
 INV_X1 _38303_ (.A(_15498_),
    .ZN(_15518_));
 INV_X1 _38304_ (.A(_15502_),
    .ZN(_15536_));
 INV_X1 _38305_ (.A(_15511_),
    .ZN(_15517_));
 INV_X1 _38306_ (.A(_15526_),
    .ZN(_15545_));
 INV_X1 _38307_ (.A(_15534_),
    .ZN(_15544_));
 INV_X1 _38308_ (.A(_15553_),
    .ZN(_15572_));
 INV_X1 _38309_ (.A(_15557_),
    .ZN(_15578_));
 INV_X1 _38310_ (.A(_15560_),
    .ZN(_15571_));
 INV_X1 _38311_ (.A(_15564_),
    .ZN(_15573_));
 INV_X1 _38312_ (.A(_15598_),
    .ZN(_15668_));
 INV_X1 _38313_ (.A(_15601_),
    .ZN(_19227_));
 INV_X1 _38314_ (.A(_15608_),
    .ZN(_15631_));
 INV_X1 _38315_ (.A(_15616_),
    .ZN(_15640_));
 INV_X1 _38316_ (.A(_15620_),
    .ZN(_15639_));
 INV_X1 _38317_ (.A(_15628_),
    .ZN(_15647_));
 INV_X1 _38318_ (.A(_15636_),
    .ZN(_15652_));
 INV_X1 _38319_ (.A(_15657_),
    .ZN(_19350_));
 INV_X1 _38320_ (.A(_15661_),
    .ZN(_19348_));
 INV_X1 _38321_ (.A(_15666_),
    .ZN(_15680_));
 INV_X1 _38322_ (.A(_15678_),
    .ZN(_19354_));
 INV_X1 _38323_ (.A(_15690_),
    .ZN(_15760_));
 INV_X1 _38324_ (.A(_15694_),
    .ZN(_15758_));
 INV_X1 _38325_ (.A(_15700_),
    .ZN(_15767_));
 INV_X1 _38326_ (.A(_15706_),
    .ZN(_19166_));
 INV_X1 _38327_ (.A(_15711_),
    .ZN(_19315_));
 INV_X1 _38328_ (.A(_15726_),
    .ZN(_15741_));
 INV_X1 _38329_ (.A(_15729_),
    .ZN(_19323_));
 INV_X1 _38330_ (.A(_15739_),
    .ZN(_15777_));
 INV_X1 _38331_ (.A(_15748_),
    .ZN(_15773_));
 INV_X1 _38332_ (.A(_15752_),
    .ZN(_15776_));
 INV_X1 _38333_ (.A(_15756_),
    .ZN(_16474_));
 INV_X1 _38334_ (.A(_15765_),
    .ZN(_16481_));
 INV_X1 _38335_ (.A(_15796_),
    .ZN(_15824_));
 INV_X1 _38336_ (.A(_15804_),
    .ZN(_15820_));
 INV_X1 _38337_ (.A(_15814_),
    .ZN(_15821_));
 INV_X1 _38338_ (.A(_15829_),
    .ZN(_15871_));
 INV_X1 _38339_ (.A(_15833_),
    .ZN(_15849_));
 INV_X1 _38340_ (.A(_15838_),
    .ZN(_15851_));
 INV_X1 _38341_ (.A(_15842_),
    .ZN(_15850_));
 INV_X1 _38342_ (.A(_15859_),
    .ZN(_15878_));
 INV_X1 _38343_ (.A(_15885_),
    .ZN(_15917_));
 INV_X1 _38344_ (.A(_15888_),
    .ZN(_15905_));
 INV_X1 _38345_ (.A(_15893_),
    .ZN(_15904_));
 INV_X1 _38346_ (.A(_15897_),
    .ZN(_15906_));
 INV_X1 _38347_ (.A(_15932_),
    .ZN(_15952_));
 INV_X1 _38348_ (.A(_15936_),
    .ZN(_15951_));
 INV_X1 _38349_ (.A(_15942_),
    .ZN(_15961_));
 INV_X1 _38350_ (.A(_15949_),
    .ZN(_15966_));
 INV_X1 _38351_ (.A(_15958_),
    .ZN(_15974_));
 INV_X1 _38352_ (.A(_15978_),
    .ZN(_19299_));
 INV_X1 _38353_ (.A(_15982_),
    .ZN(_19300_));
 INV_X1 _38354_ (.A(_15985_),
    .ZN(_19304_));
 INV_X1 _38355_ (.A(_15989_),
    .ZN(_16510_));
 INV_X1 _38356_ (.A(_15994_),
    .ZN(_16011_));
 INV_X1 _38357_ (.A(_15998_),
    .ZN(_16010_));
 INV_X1 _38358_ (.A(_16007_),
    .ZN(_16514_));
 INV_X1 _38359_ (.A(_16016_),
    .ZN(_16001_));
 INV_X1 _38360_ (.A(_16020_),
    .ZN(_16025_));
 INV_X1 _38361_ (.A(_16050_),
    .ZN(_16046_));
 INV_X1 _38362_ (.A(_16055_),
    .ZN(_16045_));
 INV_X1 _38363_ (.A(_16059_),
    .ZN(_16047_));
 INV_X1 _38364_ (.A(_16074_),
    .ZN(_16085_));
 INV_X1 _38365_ (.A(_16078_),
    .ZN(_16068_));
 INV_X1 _38366_ (.A(_16083_),
    .ZN(_16069_));
 INV_X1 _38367_ (.A(_16107_),
    .ZN(_16097_));
 INV_X1 _38368_ (.A(_16111_),
    .ZN(_16098_));
 INV_X1 _38369_ (.A(_16127_),
    .ZN(_16121_));
 INV_X1 _38370_ (.A(_16136_),
    .ZN(_16122_));
 INV_X1 _38371_ (.A(_16148_),
    .ZN(_16138_));
 INV_X1 _38372_ (.A(_16173_),
    .ZN(_16168_));
 INV_X1 _38373_ (.A(_16186_),
    .ZN(_16175_));
 INV_X1 _38374_ (.A(_16195_),
    .ZN(_16176_));
 INV_X1 _38375_ (.A(_16200_),
    .ZN(_16189_));
 INV_X1 _38376_ (.A(_16204_),
    .ZN(_19139_));
 INV_X1 _38377_ (.A(_16222_),
    .ZN(_19132_));
 INV_X1 _38378_ (.A(_16227_),
    .ZN(_19265_));
 INV_X1 _38379_ (.A(_16247_),
    .ZN(_16266_));
 INV_X1 _38380_ (.A(_16250_),
    .ZN(_19272_));
 INV_X1 _38381_ (.A(_16255_),
    .ZN(_16287_));
 INV_X1 _38382_ (.A(_16259_),
    .ZN(_16290_));
 INV_X1 _38383_ (.A(_16264_),
    .ZN(_16291_));
 INV_X1 _38384_ (.A(_16273_),
    .ZN(_16314_));
 INV_X1 _38385_ (.A(_16278_),
    .ZN(_16315_));
 INV_X1 _38386_ (.A(_16302_),
    .ZN(_16342_));
 INV_X1 _38387_ (.A(_16307_),
    .ZN(_16343_));
 INV_X1 _38388_ (.A(_16323_),
    .ZN(_16370_));
 INV_X1 _38389_ (.A(_16327_),
    .ZN(_16363_));
 INV_X1 _38390_ (.A(_16331_),
    .ZN(_16369_));
 INV_X1 _38391_ (.A(_16335_),
    .ZN(_16371_));
 INV_X1 _38392_ (.A(_16351_),
    .ZN(_16397_));
 INV_X1 _38393_ (.A(_16379_),
    .ZN(_16402_));
 INV_X1 _38394_ (.A(_16383_),
    .ZN(_16409_));
 INV_X1 _38395_ (.A(_16386_),
    .ZN(_16403_));
 INV_X1 _38396_ (.A(_16390_),
    .ZN(_16404_));
 INV_X1 _38397_ (.A(_16426_),
    .ZN(_16449_));
 INV_X1 _38398_ (.A(_16434_),
    .ZN(_16458_));
 INV_X1 _38399_ (.A(_16438_),
    .ZN(_16456_));
 INV_X1 _38400_ (.A(_16446_),
    .ZN(_16469_));
 INV_X1 _38401_ (.A(_16454_),
    .ZN(_16461_));
 INV_X1 _38402_ (.A(_16488_),
    .ZN(_19252_));
 INV_X1 _38403_ (.A(_16494_),
    .ZN(_19254_));
 INV_X1 _38404_ (.A(_16497_),
    .ZN(_19123_));
 INV_X1 _38405_ (.A(_16501_),
    .ZN(_19119_));
 INV_X1 _38406_ (.A(_16505_),
    .ZN(_19118_));
 INV_X1 _38407_ (.A(_16521_),
    .ZN(_16730_));
 INV_X1 _38408_ (.A(_16531_),
    .ZN(_16720_));
 INV_X1 _38409_ (.A(_16541_),
    .ZN(_16524_));
 INV_X1 _38410_ (.A(_16545_),
    .ZN(_19183_));
 INV_X1 _38411_ (.A(_16563_),
    .ZN(_19176_));
 INV_X1 _38412_ (.A(_16566_),
    .ZN(_18714_));
 INV_X1 _38413_ (.A(_16570_),
    .ZN(_16602_));
 INV_X1 _38414_ (.A(_16584_),
    .ZN(_16573_));
 INV_X1 _38415_ (.A(_16587_),
    .ZN(_16572_));
 INV_X1 _38416_ (.A(_16591_),
    .ZN(_16574_));
 INV_X1 _38417_ (.A(_16620_),
    .ZN(_16631_));
 INV_X1 _38418_ (.A(_16625_),
    .ZN(_16614_));
 INV_X1 _38419_ (.A(_16637_),
    .ZN(_18605_));
 INV_X1 _38420_ (.A(_16660_),
    .ZN(_17950_));
 INV_X1 _38421_ (.A(_16665_),
    .ZN(_17951_));
 INV_X1 _38422_ (.A(_16678_),
    .ZN(_16673_));
 INV_X1 _38423_ (.A(_16700_),
    .ZN(_16690_));
 INV_X1 _38424_ (.A(_16725_),
    .ZN(_19164_));
 INV_X1 _38425_ (.A(_16739_),
    .ZN(_18941_));
 INV_X1 _38426_ (.A(_16743_),
    .ZN(_18942_));
 INV_X1 _38427_ (.A(_16751_),
    .ZN(_18482_));
 INV_X1 _38428_ (.A(_16759_),
    .ZN(_16787_));
 INV_X1 _38429_ (.A(_16767_),
    .ZN(_16763_));
 INV_X1 _38430_ (.A(_16772_),
    .ZN(_16761_));
 INV_X1 _38431_ (.A(_16776_),
    .ZN(_16762_));
 INV_X1 _38432_ (.A(_16805_),
    .ZN(_16817_));
 INV_X1 _38433_ (.A(_16810_),
    .ZN(_16799_));
 INV_X1 _38434_ (.A(_16814_),
    .ZN(_16800_));
 INV_X1 _38435_ (.A(_16827_),
    .ZN(_16821_));
 INV_X1 _38436_ (.A(_16851_),
    .ZN(_16829_));
 INV_X1 _38437_ (.A(_16855_),
    .ZN(_18412_));
 INV_X1 _38438_ (.A(_16860_),
    .ZN(_16877_));
 INV_X1 _38439_ (.A(_16864_),
    .ZN(_16876_));
 INV_X1 _38440_ (.A(_16873_),
    .ZN(_18417_));
 INV_X1 _38441_ (.A(_16882_),
    .ZN(_16867_));
 INV_X1 _38442_ (.A(_16886_),
    .ZN(_16888_));
 INV_X1 _38443_ (.A(_16911_),
    .ZN(_16899_));
 INV_X1 _38444_ (.A(_16916_),
    .ZN(_16901_));
 INV_X1 _38445_ (.A(_16925_),
    .ZN(_18391_));
 INV_X1 _38446_ (.A(_16929_),
    .ZN(_18119_));
 INV_X1 _38447_ (.A(_16933_),
    .ZN(_18390_));
 INV_X1 _38448_ (.A(_16937_),
    .ZN(_18392_));
 INV_X1 _38449_ (.A(_16947_),
    .ZN(_16918_));
 INV_X1 _38450_ (.A(_16960_),
    .ZN(_18376_));
 INV_X1 _38451_ (.A(_16964_),
    .ZN(_18915_));
 INV_X1 _38452_ (.A(_16978_),
    .ZN(_18848_));
 INV_X1 _38453_ (.A(_16990_),
    .ZN(_18575_));
 INV_X1 _38454_ (.A(_16998_),
    .ZN(_17026_));
 INV_X1 _38455_ (.A(_17006_),
    .ZN(_17001_));
 INV_X1 _38456_ (.A(_17011_),
    .ZN(_17000_));
 INV_X1 _38457_ (.A(_17015_),
    .ZN(_17002_));
 INV_X1 _38458_ (.A(_17040_),
    .ZN(_17055_));
 INV_X1 _38459_ (.A(_17048_),
    .ZN(_17043_));
 INV_X1 _38460_ (.A(_17053_),
    .ZN(_17042_));
 INV_X1 _38461_ (.A(_17061_),
    .ZN(_17602_));
 INV_X1 _38462_ (.A(_17071_),
    .ZN(_17603_));
 INV_X1 _38463_ (.A(_17080_),
    .ZN(_18560_));
 INV_X1 _38464_ (.A(_17102_),
    .ZN(_17095_));
 INV_X1 _38465_ (.A(_17116_),
    .ZN(_18801_));
 INV_X1 _38466_ (.A(_17120_),
    .ZN(_18799_));
 INV_X1 _38467_ (.A(_17127_),
    .ZN(_18529_));
 INV_X1 _38468_ (.A(_17148_),
    .ZN(_17129_));
 INV_X1 _38469_ (.A(_17162_),
    .ZN(_17151_));
 INV_X1 _38470_ (.A(_17165_),
    .ZN(_17150_));
 INV_X1 _38471_ (.A(_17169_),
    .ZN(_17152_));
 INV_X1 _38472_ (.A(_17177_),
    .ZN(_17192_));
 INV_X1 _38473_ (.A(_17186_),
    .ZN(_17179_));
 INV_X1 _38474_ (.A(_17198_),
    .ZN(_18025_));
 INV_X1 _38475_ (.A(_17208_),
    .ZN(_18026_));
 INV_X1 _38476_ (.A(_17222_),
    .ZN(_17215_));
 INV_X1 _38477_ (.A(_17227_),
    .ZN(_17216_));
 INV_X1 _38478_ (.A(_17240_),
    .ZN(_17235_));
 INV_X1 _38479_ (.A(_17255_),
    .ZN(_18661_));
 INV_X1 _38480_ (.A(_17273_),
    .ZN(_17345_));
 INV_X1 _38481_ (.A(_17283_),
    .ZN(_17346_));
 INV_X1 _38482_ (.A(_17296_),
    .ZN(_17291_));
 INV_X1 _38483_ (.A(_17300_),
    .ZN(_17338_));
 INV_X1 _38484_ (.A(_17314_),
    .ZN(_17302_));
 INV_X1 _38485_ (.A(_17318_),
    .ZN(_17304_));
 INV_X1 _38486_ (.A(_17330_),
    .ZN(_17978_));
 INV_X1 _38487_ (.A(_17335_),
    .ZN(_17979_));
 INV_X1 _38488_ (.A(_17351_),
    .ZN(_18755_));
 INV_X1 _38489_ (.A(_17363_),
    .ZN(_18679_));
 INV_X1 _38490_ (.A(_17368_),
    .ZN(_18653_));
 INV_X1 _38491_ (.A(_17377_),
    .ZN(_18654_));
 INV_X1 _38492_ (.A(_17382_),
    .ZN(_17372_));
 INV_X1 _38493_ (.A(_17391_),
    .ZN(_18683_));
 INV_X1 _38494_ (.A(_17396_),
    .ZN(_17386_));
 INV_X1 _38495_ (.A(_17400_),
    .ZN(_17384_));
 INV_X1 _38496_ (.A(_17409_),
    .ZN(_17403_));
 INV_X1 _38497_ (.A(_17413_),
    .ZN(_17418_));
 INV_X1 _38498_ (.A(_17429_),
    .ZN(_18997_));
 INV_X1 _38499_ (.A(_17452_),
    .ZN(_17463_));
 INV_X1 _38500_ (.A(_17457_),
    .ZN(_17445_));
 INV_X1 _38501_ (.A(_17461_),
    .ZN(_17446_));
 INV_X1 _38502_ (.A(_17473_),
    .ZN(_17858_));
 INV_X1 _38503_ (.A(_17477_),
    .ZN(_17843_));
 INV_X1 _38504_ (.A(_17480_),
    .ZN(_17859_));
 INV_X1 _38505_ (.A(_17484_),
    .ZN(_17857_));
 INV_X1 _38506_ (.A(_17498_),
    .ZN(_17491_));
 INV_X1 _38507_ (.A(_17506_),
    .ZN(_17493_));
 INV_X1 _38508_ (.A(_17520_),
    .ZN(_17509_));
 INV_X1 _38509_ (.A(_17524_),
    .ZN(_17510_));
 INV_X1 _38510_ (.A(_17541_),
    .ZN(_17536_));
 INV_X1 _38511_ (.A(_17550_),
    .ZN(_17535_));
 INV_X1 _38512_ (.A(_17560_),
    .ZN(_17552_));
 INV_X1 _38513_ (.A(_17574_),
    .ZN(_17562_));
 INV_X1 _38514_ (.A(_17587_),
    .ZN(_17580_));
 INV_X1 _38515_ (.A(_17592_),
    .ZN(_17581_));
 INV_X1 _38516_ (.A(_17596_),
    .ZN(_17582_));
 INV_X1 _38517_ (.A(_17607_),
    .ZN(_18525_));
 INV_X1 _38518_ (.A(_17612_),
    .ZN(_17625_));
 INV_X1 _38519_ (.A(_17616_),
    .ZN(_17623_));
 INV_X1 _38520_ (.A(_17628_),
    .ZN(_17619_));
 INV_X1 _38521_ (.A(_17646_),
    .ZN(_17654_));
 INV_X1 _38522_ (.A(_17659_),
    .ZN(_17648_));
 INV_X1 _38523_ (.A(_17664_),
    .ZN(_18632_));
 INV_X1 _38524_ (.A(_17668_),
    .ZN(_18631_));
 INV_X1 _38525_ (.A(_17673_),
    .ZN(_19028_));
 INV_X1 _38526_ (.A(_17685_),
    .ZN(_18362_));
 INV_X1 _38527_ (.A(_17710_),
    .ZN(_17692_));
 INV_X1 _38528_ (.A(_17718_),
    .ZN(_17712_));
 INV_X1 _38529_ (.A(_17723_),
    .ZN(_17713_));
 INV_X1 _38530_ (.A(_17727_),
    .ZN(_17714_));
 INV_X1 _38531_ (.A(_17739_),
    .ZN(_17750_));
 INV_X1 _38532_ (.A(_17743_),
    .ZN(_17733_));
 INV_X1 _38533_ (.A(_17748_),
    .ZN(_17734_));
 INV_X1 _38534_ (.A(_17764_),
    .ZN(_17757_));
 INV_X1 _38535_ (.A(_17769_),
    .ZN(_17758_));
 INV_X1 _38536_ (.A(_17773_),
    .ZN(_17759_));
 INV_X1 _38537_ (.A(_17786_),
    .ZN(_17781_));
 INV_X1 _38538_ (.A(_17795_),
    .ZN(_17779_));
 INV_X1 _38539_ (.A(_17800_),
    .ZN(_18218_));
 INV_X1 _38540_ (.A(_17804_),
    .ZN(_18339_));
 INV_X1 _38541_ (.A(_17809_),
    .ZN(_18338_));
 INV_X1 _38542_ (.A(_17819_),
    .ZN(_17811_));
 INV_X1 _38543_ (.A(_17822_),
    .ZN(_18988_));
 INV_X1 _38544_ (.A(_17827_),
    .ZN(_18308_));
 INV_X1 _38545_ (.A(_17831_),
    .ZN(_18306_));
 INV_X1 _38546_ (.A(_17840_),
    .ZN(_18310_));
 INV_X1 _38547_ (.A(_17873_),
    .ZN(_17861_));
 INV_X1 _38548_ (.A(_17878_),
    .ZN(_17863_));
 INV_X1 _38549_ (.A(_17891_),
    .ZN(_17881_));
 INV_X1 _38550_ (.A(_17909_),
    .ZN(_17903_));
 INV_X1 _38551_ (.A(_17923_),
    .ZN(_17911_));
 INV_X1 _38552_ (.A(_17933_),
    .ZN(_17925_));
 INV_X1 _38553_ (.A(_17941_),
    .ZN(_17927_));
 INV_X1 _38554_ (.A(_17959_),
    .ZN(_17954_));
 INV_X1 _38555_ (.A(_17964_),
    .ZN(_17953_));
 INV_X1 _38556_ (.A(_17968_),
    .ZN(_17955_));
 INV_X1 _38557_ (.A(_17983_),
    .ZN(_18503_));
 INV_X1 _38558_ (.A(_17988_),
    .ZN(_18504_));
 INV_X1 _38559_ (.A(_17998_),
    .ZN(_17990_));
 INV_X1 _38560_ (.A(_18011_),
    .ZN(_18003_));
 INV_X1 _38561_ (.A(_18015_),
    .ZN(_18004_));
 INV_X1 _38562_ (.A(_18019_),
    .ZN(_18005_));
 INV_X1 _38563_ (.A(_18030_),
    .ZN(_18553_));
 INV_X1 _38564_ (.A(_18035_),
    .ZN(_18552_));
 INV_X1 _38565_ (.A(_18045_),
    .ZN(_18038_));
 INV_X1 _38566_ (.A(_18054_),
    .ZN(_18579_));
 INV_X1 _38567_ (.A(_18059_),
    .ZN(_18047_));
 INV_X1 _38568_ (.A(_18063_),
    .ZN(_18048_));
 INV_X1 _38569_ (.A(_18070_),
    .ZN(_18066_));
 INV_X1 _38570_ (.A(_18075_),
    .ZN(_18907_));
 INV_X1 _38571_ (.A(_18089_),
    .ZN(_18082_));
 INV_X1 _38572_ (.A(_18092_),
    .ZN(_18081_));
 INV_X1 _38573_ (.A(_18096_),
    .ZN(_18083_));
 INV_X1 _38574_ (.A(_18113_),
    .ZN(_18106_));
 INV_X1 _38575_ (.A(_18134_),
    .ZN(_18478_));
 INV_X1 _38576_ (.A(_18139_),
    .ZN(_18152_));
 INV_X1 _38577_ (.A(_18143_),
    .ZN(_18151_));
 INV_X1 _38578_ (.A(_18155_),
    .ZN(_18146_));
 INV_X1 _38579_ (.A(_18160_),
    .ZN(_18282_));
 INV_X1 _38580_ (.A(_18164_),
    .ZN(_19003_));
 INV_X1 _38581_ (.A(_18185_),
    .ZN(_18176_));
 INV_X1 _38582_ (.A(_18194_),
    .ZN(_18187_));
 INV_X1 _38583_ (.A(_18203_),
    .ZN(_18346_));
 INV_X1 _38584_ (.A(_18225_),
    .ZN(_18597_));
 INV_X1 _38585_ (.A(_18234_),
    .ZN(_18598_));
 INV_X1 _38586_ (.A(_18239_),
    .ZN(_18227_));
 INV_X1 _38587_ (.A(_18243_),
    .ZN(_18895_));
 INV_X1 _38588_ (.A(_18247_),
    .ZN(_18894_));
 INV_X1 _38589_ (.A(_18259_),
    .ZN(_18365_));
 INV_X1 _38590_ (.A(_18264_),
    .ZN(_18254_));
 INV_X1 _38591_ (.A(_18268_),
    .ZN(_18252_));
 INV_X1 _38592_ (.A(_18275_),
    .ZN(_18271_));
 INV_X1 _38593_ (.A(_18317_),
    .ZN(_18986_));
 INV_X1 _38594_ (.A(_18325_),
    .ZN(_19039_));
 INV_X1 _38595_ (.A(_18332_),
    .ZN(_19045_));
 INV_X1 _38596_ (.A(_18369_),
    .ZN(_19030_));
 INV_X1 _38597_ (.A(_18382_),
    .ZN(_17563_));
 INV_X1 _38598_ (.A(_18421_),
    .ZN(_18899_));
 INV_X1 _38599_ (.A(_18426_),
    .ZN(_18955_));
 INV_X1 _38600_ (.A(_18431_),
    .ZN(_18442_));
 INV_X1 _38601_ (.A(_18434_),
    .ZN(_18961_));
 INV_X1 _38602_ (.A(_18450_),
    .ZN(_18459_));
 INV_X1 _38603_ (.A(_18485_),
    .ZN(_18946_));
 INV_X1 _38604_ (.A(_18490_),
    .ZN(_18815_));
 INV_X1 _38605_ (.A(_18497_),
    .ZN(_18823_));
 INV_X1 _38606_ (.A(_18534_),
    .ZN(_18806_));
 INV_X1 _38607_ (.A(_18539_),
    .ZN(_18859_));
 INV_X1 _38608_ (.A(_18546_),
    .ZN(_18868_));
 INV_X1 _38609_ (.A(_18583_),
    .ZN(_18851_));
 INV_X1 _38610_ (.A(_18588_),
    .ZN(_18723_));
 INV_X1 _38611_ (.A(_18591_),
    .ZN(_18730_));
 INV_X1 _38612_ (.A(_18617_),
    .ZN(_18627_));
 INV_X1 _38613_ (.A(_18635_),
    .ZN(_18709_));
 INV_X1 _38614_ (.A(_18639_),
    .ZN(_18707_));
 INV_X1 _38615_ (.A(_18644_),
    .ZN(_18766_));
 INV_X1 _38616_ (.A(_18647_),
    .ZN(_18774_));
 INV_X1 _38617_ (.A(_18687_),
    .ZN(_18758_));
 INV_X1 _38618_ (.A(_18689_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[11] ));
 INV_X1 _38619_ (.A(_18691_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[12] ));
 INV_X1 _38620_ (.A(_18693_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[13] ));
 INV_X1 _38621_ (.A(_18695_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[14] ));
 INV_X1 _38622_ (.A(_18697_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[15] ));
 INV_X1 _38623_ (.A(_18699_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[16] ));
 INV_X1 _38624_ (.A(_18701_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[17] ));
 INV_X1 _38625_ (.A(_18705_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[18] ));
 INV_X1 _38626_ (.A(_18710_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[19] ));
 INV_X1 _38627_ (.A(_18715_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[20] ));
 INV_X1 _38628_ (.A(_18724_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[6] ));
 INV_X1 _38629_ (.A(_18727_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[7] ));
 INV_X1 _38630_ (.A(_18731_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[8] ));
 INV_X1 _38631_ (.A(_18733_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[9] ));
 INV_X1 _38632_ (.A(_18735_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[10] ));
 INV_X1 _38633_ (.A(_18737_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[11] ));
 INV_X1 _38634_ (.A(_18739_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[12] ));
 INV_X1 _38635_ (.A(_18741_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[13] ));
 INV_X1 _38636_ (.A(_18743_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[14] ));
 INV_X1 _38637_ (.A(_18745_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[15] ));
 INV_X1 _38638_ (.A(_18747_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[16] ));
 INV_X1 _38639_ (.A(_18749_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[17] ));
 INV_X1 _38640_ (.A(_18753_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[18] ));
 INV_X1 _38641_ (.A(_18759_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[20] ));
 INV_X1 _38642_ (.A(_18768_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[6] ));
 INV_X1 _38643_ (.A(_18771_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[7] ));
 INV_X1 _38644_ (.A(_18775_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[8] ));
 INV_X1 _38645_ (.A(_18777_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[9] ));
 INV_X1 _38646_ (.A(_18779_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[10] ));
 INV_X1 _38647_ (.A(_18781_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[11] ));
 INV_X1 _38648_ (.A(_18783_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[12] ));
 INV_X1 _38649_ (.A(_18785_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[13] ));
 INV_X1 _38650_ (.A(_18787_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[14] ));
 INV_X1 _38651_ (.A(_18789_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[15] ));
 INV_X1 _38652_ (.A(_18791_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[16] ));
 INV_X1 _38653_ (.A(_18793_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[17] ));
 INV_X1 _38654_ (.A(_18797_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[18] ));
 INV_X1 _38655_ (.A(_18802_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[19] ));
 INV_X1 _38656_ (.A(_18807_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[20] ));
 INV_X1 _38657_ (.A(_18816_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[6] ));
 INV_X1 _38658_ (.A(_18820_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[7] ));
 INV_X1 _38659_ (.A(_18824_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[8] ));
 INV_X1 _38660_ (.A(_18826_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[9] ));
 INV_X1 _38661_ (.A(_18828_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[10] ));
 INV_X1 _38662_ (.A(_18830_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[11] ));
 INV_X1 _38663_ (.A(_18832_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[12] ));
 INV_X1 _38664_ (.A(_18834_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[13] ));
 INV_X1 _38665_ (.A(_18836_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[14] ));
 INV_X1 _38666_ (.A(_18838_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[15] ));
 INV_X1 _38667_ (.A(_18840_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[16] ));
 INV_X1 _38668_ (.A(_18842_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[17] ));
 INV_X1 _38669_ (.A(_18846_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[18] ));
 INV_X1 _38670_ (.A(_18852_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[20] ));
 INV_X1 _38671_ (.A(_18861_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[6] ));
 INV_X1 _38672_ (.A(_18865_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[7] ));
 INV_X1 _38673_ (.A(_18869_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[8] ));
 INV_X1 _38674_ (.A(_18871_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[9] ));
 INV_X1 _38675_ (.A(_18873_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[10] ));
 INV_X1 _38676_ (.A(_18875_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[11] ));
 INV_X1 _38677_ (.A(_18877_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[12] ));
 INV_X1 _38678_ (.A(_18879_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[13] ));
 INV_X1 _38679_ (.A(_18881_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[14] ));
 INV_X1 _38680_ (.A(_18883_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[15] ));
 INV_X1 _38681_ (.A(_18885_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[16] ));
 INV_X1 _38682_ (.A(_18887_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[17] ));
 INV_X1 _38683_ (.A(_18891_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[18] ));
 INV_X1 _38684_ (.A(_18896_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[19] ));
 INV_X1 _38685_ (.A(_18900_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[20] ));
 INV_X1 _38686_ (.A(_18909_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[6] ));
 INV_X1 _38687_ (.A(_18912_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[7] ));
 INV_X1 _38688_ (.A(_18916_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[8] ));
 INV_X1 _38689_ (.A(_18918_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[9] ));
 INV_X1 _38690_ (.A(_18920_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[10] ));
 INV_X1 _38691_ (.A(_18922_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[11] ));
 INV_X1 _38692_ (.A(_18924_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[12] ));
 INV_X1 _38693_ (.A(_18926_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[13] ));
 INV_X1 _38694_ (.A(_18928_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[14] ));
 INV_X1 _38695_ (.A(_18930_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[15] ));
 INV_X1 _38696_ (.A(_18932_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[16] ));
 INV_X1 _38697_ (.A(_18934_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[17] ));
 INV_X1 _38698_ (.A(_18938_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[18] ));
 INV_X1 _38699_ (.A(_18943_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[19] ));
 INV_X1 _38700_ (.A(_18947_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[20] ));
 INV_X1 _38701_ (.A(_18956_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[6] ));
 INV_X1 _38702_ (.A(_18959_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[7] ));
 INV_X1 _38703_ (.A(_18962_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[8] ));
 INV_X1 _38704_ (.A(_18964_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[9] ));
 INV_X1 _38705_ (.A(_18966_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[10] ));
 INV_X1 _38706_ (.A(_18968_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[11] ));
 INV_X1 _38707_ (.A(_18970_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[12] ));
 INV_X1 _38708_ (.A(_18972_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[13] ));
 INV_X1 _38709_ (.A(_18974_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[14] ));
 INV_X1 _38710_ (.A(_18976_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[15] ));
 INV_X1 _38711_ (.A(_18978_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[16] ));
 INV_X1 _38712_ (.A(_18980_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[17] ));
 INV_X1 _38713_ (.A(_18984_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[18] ));
 INV_X1 _38714_ (.A(_18989_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[20] ));
 INV_X1 _38715_ (.A(_18998_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[6] ));
 INV_X1 _38716_ (.A(_19001_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[7] ));
 INV_X1 _38717_ (.A(_19004_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[8] ));
 INV_X1 _38718_ (.A(_19006_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[9] ));
 INV_X1 _38719_ (.A(_19008_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[10] ));
 INV_X1 _38720_ (.A(_19010_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[11] ));
 INV_X1 _38721_ (.A(_19012_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[12] ));
 INV_X1 _38722_ (.A(_19014_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[13] ));
 INV_X1 _38723_ (.A(_19016_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[14] ));
 INV_X1 _38724_ (.A(_19018_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[15] ));
 INV_X1 _38725_ (.A(_19020_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[16] ));
 INV_X1 _38726_ (.A(_19022_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[17] ));
 INV_X1 _38727_ (.A(_19026_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[18] ));
 INV_X1 _38728_ (.A(_19031_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[20] ));
 INV_X1 _38729_ (.A(_19040_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[6] ));
 INV_X1 _38730_ (.A(_19043_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[7] ));
 INV_X1 _38731_ (.A(_19047_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[8] ));
 INV_X1 _38732_ (.A(_19049_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[9] ));
 INV_X1 _38733_ (.A(_19051_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[10] ));
 INV_X1 _38734_ (.A(_19053_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[11] ));
 INV_X1 _38735_ (.A(_19055_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[12] ));
 INV_X1 _38736_ (.A(_19057_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[13] ));
 INV_X1 _38737_ (.A(_19059_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[14] ));
 INV_X1 _38738_ (.A(_19061_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[15] ));
 INV_X1 _38739_ (.A(_19063_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[16] ));
 INV_X1 _38740_ (.A(_19065_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[17] ));
 INV_X1 _38741_ (.A(_19069_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[18] ));
 INV_X1 _38742_ (.A(_19074_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[20] ));
 INV_X1 _38743_ (.A(_19079_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[4] ));
 INV_X1 _38744_ (.A(_19085_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[6] ));
 INV_X1 _38745_ (.A(_19089_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[7] ));
 INV_X1 _38746_ (.A(_19093_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[8] ));
 INV_X1 _38747_ (.A(_19095_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[9] ));
 INV_X1 _38748_ (.A(_19097_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[10] ));
 INV_X1 _38749_ (.A(_19099_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[11] ));
 INV_X1 _38750_ (.A(_19101_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[12] ));
 INV_X1 _38751_ (.A(_19103_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[13] ));
 INV_X1 _38752_ (.A(_19105_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[14] ));
 INV_X1 _38753_ (.A(_19107_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[15] ));
 INV_X1 _38754_ (.A(_19109_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[16] ));
 INV_X1 _38755_ (.A(_19111_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[17] ));
 INV_X1 _38756_ (.A(_19115_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[18] ));
 INV_X1 _38757_ (.A(_19120_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[19] ));
 INV_X1 _38758_ (.A(_19124_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[20] ));
 INV_X1 _38759_ (.A(_19133_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[6] ));
 INV_X1 _38760_ (.A(_19136_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[7] ));
 INV_X1 _38761_ (.A(_19140_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[8] ));
 INV_X1 _38762_ (.A(_19142_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[9] ));
 INV_X1 _38763_ (.A(_19144_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[10] ));
 INV_X1 _38764_ (.A(_19146_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[11] ));
 INV_X1 _38765_ (.A(_19148_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[12] ));
 INV_X1 _38766_ (.A(_19150_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[13] ));
 INV_X1 _38767_ (.A(_19152_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[14] ));
 INV_X1 _38768_ (.A(_19154_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[15] ));
 INV_X1 _38769_ (.A(_19156_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[16] ));
 INV_X1 _38770_ (.A(_19158_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[17] ));
 INV_X1 _38771_ (.A(_19162_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[18] ));
 INV_X1 _38772_ (.A(_19167_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[20] ));
 INV_X1 _38773_ (.A(_19172_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[4] ));
 INV_X1 _38774_ (.A(_19178_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[6] ));
 INV_X1 _38775_ (.A(_19181_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[7] ));
 INV_X1 _38776_ (.A(_19184_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[8] ));
 INV_X1 _38777_ (.A(_19186_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[9] ));
 INV_X1 _38778_ (.A(_19188_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[10] ));
 INV_X1 _38779_ (.A(_19190_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[11] ));
 INV_X1 _38780_ (.A(_19192_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[12] ));
 INV_X1 _38781_ (.A(_19194_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[13] ));
 INV_X1 _38782_ (.A(_19196_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[14] ));
 INV_X1 _38783_ (.A(_19198_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[15] ));
 INV_X1 _38784_ (.A(_19200_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[16] ));
 INV_X1 _38785_ (.A(_19202_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[17] ));
 INV_X1 _38786_ (.A(_19206_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[18] ));
 INV_X1 _38787_ (.A(_19211_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[20] ));
 INV_X1 _38788_ (.A(_19216_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[4] ));
 INV_X1 _38789_ (.A(_19222_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[6] ));
 INV_X1 _38790_ (.A(_19225_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[7] ));
 INV_X1 _38791_ (.A(_19228_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[8] ));
 INV_X1 _38792_ (.A(_19230_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[9] ));
 INV_X1 _38793_ (.A(_19232_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[10] ));
 INV_X1 _38794_ (.A(_19234_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[11] ));
 INV_X1 _38795_ (.A(_19236_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[12] ));
 INV_X1 _38796_ (.A(_19238_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[13] ));
 INV_X1 _38797_ (.A(_19240_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[14] ));
 INV_X1 _38798_ (.A(_19242_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[15] ));
 INV_X1 _38799_ (.A(_19244_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[16] ));
 INV_X1 _38800_ (.A(_19246_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[17] ));
 INV_X1 _38801_ (.A(_19250_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[18] ));
 INV_X1 _38802_ (.A(_19255_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[20] ));
 INV_X1 _38803_ (.A(_19260_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[4] ));
 INV_X1 _38804_ (.A(_19266_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[6] ));
 INV_X1 _38805_ (.A(_19270_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[7] ));
 INV_X1 _38806_ (.A(_19274_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[8] ));
 INV_X1 _38807_ (.A(_19276_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[9] ));
 INV_X1 _38808_ (.A(_19278_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[10] ));
 INV_X1 _38809_ (.A(_19280_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[11] ));
 INV_X1 _38810_ (.A(_19282_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[12] ));
 INV_X1 _38811_ (.A(_19284_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[13] ));
 INV_X1 _38812_ (.A(_19286_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[14] ));
 INV_X1 _38813_ (.A(_19288_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[15] ));
 INV_X1 _38814_ (.A(_19290_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[16] ));
 INV_X1 _38815_ (.A(_19292_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[17] ));
 INV_X1 _38816_ (.A(_19296_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[18] ));
 INV_X1 _38817_ (.A(_19301_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[19] ));
 INV_X1 _38818_ (.A(_19305_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[20] ));
 INV_X1 _38819_ (.A(_19310_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[4] ));
 INV_X1 _38820_ (.A(_19316_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[6] ));
 INV_X1 _38821_ (.A(_19320_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[7] ));
 INV_X1 _38822_ (.A(_19324_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[8] ));
 INV_X1 _38823_ (.A(_19326_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[9] ));
 INV_X1 _38824_ (.A(_19328_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[10] ));
 INV_X1 _38825_ (.A(_19330_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[11] ));
 INV_X1 _38826_ (.A(_19332_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[12] ));
 INV_X1 _38827_ (.A(_19334_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[13] ));
 INV_X1 _38828_ (.A(_19336_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[14] ));
 INV_X1 _38829_ (.A(_19338_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[15] ));
 INV_X1 _38830_ (.A(_19340_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[16] ));
 INV_X1 _38831_ (.A(_19342_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[17] ));
 INV_X1 _38832_ (.A(_19346_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[18] ));
 INV_X1 _38833_ (.A(_19351_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[19] ));
 INV_X1 _38834_ (.A(_19355_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[20] ));
 INV_X1 _38835_ (.A(_19360_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[4] ));
 INV_X1 _38836_ (.A(_19366_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[6] ));
 INV_X1 _38837_ (.A(_19369_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[7] ));
 INV_X1 _38838_ (.A(_19372_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[8] ));
 INV_X1 _38839_ (.A(_19374_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[9] ));
 INV_X1 _38840_ (.A(_19376_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[10] ));
 INV_X1 _38841_ (.A(_19378_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[11] ));
 INV_X1 _38842_ (.A(_19380_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[12] ));
 INV_X1 _38843_ (.A(_19382_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[13] ));
 INV_X1 _38844_ (.A(_19384_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[14] ));
 INV_X1 _38845_ (.A(_19386_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[15] ));
 INV_X1 _38846_ (.A(_19388_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[16] ));
 INV_X1 _38847_ (.A(_19390_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[17] ));
 INV_X1 _38848_ (.A(_19394_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[18] ));
 INV_X1 _38849_ (.A(_19399_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[20] ));
 INV_X1 _38850_ (.A(_19404_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[4] ));
 INV_X1 _38851_ (.A(_19410_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[6] ));
 INV_X1 _38852_ (.A(_19414_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[7] ));
 INV_X1 _38853_ (.A(_19418_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[8] ));
 INV_X1 _38854_ (.A(_19420_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[9] ));
 INV_X1 _38855_ (.A(_19422_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[10] ));
 INV_X1 _38856_ (.A(_06747_),
    .ZN(_19433_));
 INV_X1 _38857_ (.A(_06759_),
    .ZN(_19437_));
 INV_X1 _38858_ (.A(_14219_),
    .ZN(_19481_));
 INV_X1 _38859_ (.A(_14238_),
    .ZN(_19538_));
 INV_X1 _38860_ (.A(_14257_),
    .ZN(_19595_));
 INV_X1 _38861_ (.A(_14282_),
    .ZN(_19652_));
 INV_X1 _38862_ (.A(_14281_),
    .ZN(_19658_));
 INV_X1 _38863_ (.A(_07494_),
    .ZN(_19665_));
 INV_X1 _38864_ (.A(_14299_),
    .ZN(_19709_));
 INV_X1 _38865_ (.A(_14298_),
    .ZN(_19715_));
 INV_X1 _38866_ (.A(_14316_),
    .ZN(_19766_));
 INV_X1 _38867_ (.A(_14315_),
    .ZN(_19772_));
 INV_X1 _38868_ (.A(_14328_),
    .ZN(_19823_));
 INV_X1 _38869_ (.A(_14345_),
    .ZN(_19880_));
 INV_X1 _38870_ (.A(_14349_),
    .ZN(_19886_));
 INV_X1 _38871_ (.A(_14367_),
    .ZN(_19937_));
 INV_X1 _38872_ (.A(_14366_),
    .ZN(_19943_));
 INV_X1 _38873_ (.A(_14379_),
    .ZN(_19994_));
 INV_X1 _38874_ (.A(_14401_),
    .ZN(_20051_));
 INV_X1 _38875_ (.A(_14400_),
    .ZN(_20057_));
 INV_X1 _38876_ (.A(_14413_),
    .ZN(_20108_));
 INV_X1 _38877_ (.A(_14435_),
    .ZN(_20165_));
 INV_X1 _38878_ (.A(_14452_),
    .ZN(_20222_));
 INV_X1 _38879_ (.A(_14451_),
    .ZN(_20228_));
 INV_X1 _38880_ (.A(_14464_),
    .ZN(_20279_));
 INV_X1 _38881_ (.A(_14481_),
    .ZN(_20336_));
 AND2_X1 _38882_ (.A1(_00448_),
    .A2(_10394_),
    .ZN(_11980_));
 BUF_X4 _38883_ (.A(_10268_),
    .Z(_11981_));
 AOI21_X4 _38884_ (.A(_11980_),
    .B1(_11981_),
    .B2(_20386_),
    .ZN(_14493_));
 AND2_X1 _38885_ (.A1(_00460_),
    .A2(_10394_),
    .ZN(_11982_));
 AOI21_X2 _38886_ (.A(_11982_),
    .B1(_11981_),
    .B2(_20365_),
    .ZN(_20409_));
 AND2_X1 _38887_ (.A1(_20371_),
    .A2(_11981_),
    .ZN(_11983_));
 AOI21_X2 _38888_ (.A(_11983_),
    .B1(_10394_),
    .B2(_00457_),
    .ZN(_20423_));
 AND2_X1 _38889_ (.A1(_20377_),
    .A2(_11981_),
    .ZN(_11984_));
 AOI21_X2 _38890_ (.A(_11984_),
    .B1(_10394_),
    .B2(_00455_),
    .ZN(_20437_));
 AND2_X1 _38891_ (.A1(_00452_),
    .A2(_10394_),
    .ZN(_11985_));
 AOI21_X2 _38892_ (.A(_11985_),
    .B1(_11981_),
    .B2(_20383_),
    .ZN(_20406_));
 AND2_X1 _38893_ (.A1(_20389_),
    .A2(_10394_),
    .ZN(_11986_));
 AOI21_X2 _38894_ (.A(_11986_),
    .B1(_11981_),
    .B2(_00449_),
    .ZN(_20462_));
 NOR2_X1 _38895_ (.A1(_10617_),
    .A2(_10665_),
    .ZN(_11987_));
 OAI21_X2 _38896_ (.A(_10795_),
    .B1(_10657_),
    .B2(_11987_),
    .ZN(_20466_));
 INV_X1 _38897_ (.A(_14500_),
    .ZN(_14505_));
 INV_X1 _38898_ (.A(_10934_),
    .ZN(_20492_));
 INV_X1 _38899_ (.A(_10941_),
    .ZN(_20496_));
 BUF_X2 _38900_ (.A(_11060_),
    .Z(_11988_));
 NOR2_X1 _38901_ (.A1(_11099_),
    .A2(_11988_),
    .ZN(_11989_));
 AOI21_X2 _38902_ (.A(_11989_),
    .B1(_11988_),
    .B2(_00468_),
    .ZN(_20574_));
 AND2_X1 _38903_ (.A1(_00470_),
    .A2(_11988_),
    .ZN(_11990_));
 BUF_X4 _38904_ (.A(_11012_),
    .Z(_11991_));
 AOI21_X2 _38905_ (.A(_11990_),
    .B1(_11991_),
    .B2(_20518_),
    .ZN(_20588_));
 AND2_X1 _38906_ (.A1(_00466_),
    .A2(_11988_),
    .ZN(_11992_));
 AOI21_X2 _38907_ (.A(_11992_),
    .B1(_11991_),
    .B2(_20533_),
    .ZN(_20549_));
 NOR2_X1 _38908_ (.A1(_11110_),
    .A2(_11988_),
    .ZN(_11993_));
 AOI21_X2 _38909_ (.A(_11993_),
    .B1(_11988_),
    .B2(_00465_),
    .ZN(_20598_));
 AND2_X1 _38910_ (.A1(_00463_),
    .A2(_11988_),
    .ZN(_11994_));
 AOI21_X2 _38911_ (.A(_11994_),
    .B1(_11991_),
    .B2(_00464_),
    .ZN(_20606_));
 NAND2_X2 _38912_ (.A1(_11314_),
    .A2(_11351_),
    .ZN(_20610_));
 INV_X1 _38913_ (.A(_11526_),
    .ZN(_20624_));
 INV_X1 _38914_ (.A(_11613_),
    .ZN(_20640_));
 AND2_X1 _38915_ (.A1(_11684_),
    .A2(_11755_),
    .ZN(_20762_));
 INV_X1 _38916_ (.A(_16475_),
    .ZN(_16727_));
 AND2_X1 _38917_ (.A1(_11825_),
    .A2(_11844_),
    .ZN(_20800_));
 AND2_X1 _38918_ (.A1(_11654_),
    .A2(_11882_),
    .ZN(_20871_));
 AND2_X1 _38919_ (.A1(_11643_),
    .A2(_11685_),
    .ZN(_20879_));
 BUF_X1 _38920_ (.A(_12193_),
    .Z(_11995_));
 MUX2_X1 _38921_ (.A(_12216_),
    .B(_12209_),
    .S(_11995_),
    .Z(_21157_));
 MUX2_X1 _38922_ (.A(_00476_),
    .B(_21154_),
    .S(_11995_),
    .Z(_11996_));
 INV_X2 _38923_ (.A(_11996_),
    .ZN(_14060_));
 MUX2_X1 _38924_ (.A(_00488_),
    .B(_21133_),
    .S(_11995_),
    .Z(_11997_));
 INV_X1 _38925_ (.A(_11997_),
    .ZN(_21171_));
 MUX2_X1 _38926_ (.A(_00482_),
    .B(_21142_),
    .S(_11995_),
    .Z(_11998_));
 INV_X1 _38927_ (.A(_11998_),
    .ZN(_21192_));
 MUX2_X1 _38928_ (.A(_00483_),
    .B(_21145_),
    .S(_11995_),
    .Z(_11999_));
 INV_X1 _38929_ (.A(_11999_),
    .ZN(_21199_));
 MUX2_X1 _38930_ (.A(_00479_),
    .B(_21148_),
    .S(_11995_),
    .Z(_12000_));
 INV_X1 _38931_ (.A(_12000_),
    .ZN(_21216_));
 MUX2_X1 _38932_ (.A(_00477_),
    .B(_00478_),
    .S(_11995_),
    .Z(_12001_));
 INV_X1 _38933_ (.A(_12001_),
    .ZN(_21224_));
 AND3_X1 _38934_ (.A1(_12433_),
    .A2(_12455_),
    .A3(_12542_),
    .ZN(_12002_));
 OAI21_X2 _38935_ (.A(_12644_),
    .B1(_12002_),
    .B2(_12501_),
    .ZN(_21228_));
 INV_X1 _38936_ (.A(_12800_),
    .ZN(_14067_));
 INV_X1 _38937_ (.A(_12792_),
    .ZN(_21254_));
 AND2_X1 _38938_ (.A1(_00490_),
    .A2(_12877_),
    .ZN(_12003_));
 BUF_X4 _38939_ (.A(_13180_),
    .Z(_12004_));
 AOI21_X4 _38940_ (.A(_12003_),
    .B1(_12004_),
    .B2(_21295_),
    .ZN(_14075_));
 MUX2_X1 _38941_ (.A(_13003_),
    .B(_13004_),
    .S(_12004_),
    .Z(_21315_));
 AND2_X1 _38942_ (.A1(_00491_),
    .A2(_13180_),
    .ZN(_12005_));
 AOI21_X2 _38943_ (.A(_12005_),
    .B1(_12877_),
    .B2(_21298_),
    .ZN(_21371_));
 INV_X1 _38944_ (.A(_00843_),
    .ZN(_21389_));
 INV_X1 _38945_ (.A(_00918_),
    .ZN(_14082_));
 INV_X1 _38946_ (.A(_00678_),
    .ZN(_21405_));
 BUF_X1 _38947_ (.A(_00995_),
    .Z(_12006_));
 AND2_X1 _38948_ (.A1(_21442_),
    .A2(_12006_),
    .ZN(_12007_));
 AOI21_X4 _38949_ (.A(_12007_),
    .B1(_01104_),
    .B2(_00504_),
    .ZN(_14090_));
 MUX2_X1 _38950_ (.A(_00508_),
    .B(_21439_),
    .S(_12006_),
    .Z(_12008_));
 INV_X1 _38951_ (.A(_12008_),
    .ZN(_21462_));
 MUX2_X1 _38952_ (.A(_21445_),
    .B(_00505_),
    .S(_12006_),
    .Z(_12009_));
 INV_X1 _38953_ (.A(_12009_),
    .ZN(_21518_));
 NAND2_X2 _38954_ (.A1(_01597_),
    .A2(_01529_),
    .ZN(_21522_));
 INV_X1 _38955_ (.A(_01614_),
    .ZN(_21530_));
 INV_X1 _38956_ (.A(_01732_),
    .ZN(_14097_));
 INV_X1 _38957_ (.A(_01724_),
    .ZN(_21548_));
 INV_X1 _38958_ (.A(_01731_),
    .ZN(_21552_));
 BUF_X1 _38959_ (.A(_01805_),
    .Z(_12010_));
 MUX2_X1 _38960_ (.A(_01874_),
    .B(_01868_),
    .S(_12010_),
    .Z(_21595_));
 MUX2_X1 _38961_ (.A(_00518_),
    .B(_21592_),
    .S(_12010_),
    .Z(_12011_));
 INV_X2 _38962_ (.A(_12011_),
    .ZN(_14105_));
 MUX2_X1 _38963_ (.A(_00521_),
    .B(_21586_),
    .S(_12010_),
    .Z(_12012_));
 INV_X1 _38964_ (.A(_12012_),
    .ZN(_21654_));
 MUX2_X1 _38965_ (.A(_00519_),
    .B(_00520_),
    .S(_12010_),
    .Z(_12013_));
 INV_X1 _38966_ (.A(_12013_),
    .ZN(_21662_));
 CLKBUF_X3 _38967_ (.A(_02533_),
    .Z(_12014_));
 MUX2_X1 _38968_ (.A(_21733_),
    .B(_00532_),
    .S(_12014_),
    .Z(_12015_));
 INV_X2 _38969_ (.A(_12015_),
    .ZN(_14120_));
 MUX2_X1 _38970_ (.A(_21730_),
    .B(_00536_),
    .S(_12014_),
    .Z(_12016_));
 INV_X1 _38971_ (.A(_12016_),
    .ZN(_21753_));
 MUX2_X1 _38972_ (.A(_00533_),
    .B(_21736_),
    .S(_12014_),
    .Z(_12017_));
 INV_X1 _38973_ (.A(_12017_),
    .ZN(_21809_));
 NAND2_X1 _38974_ (.A1(_02838_),
    .A2(_03008_),
    .ZN(_12018_));
 OAI21_X1 _38975_ (.A(_02765_),
    .B1(_12018_),
    .B2(_03018_),
    .ZN(_12019_));
 OAI21_X2 _38976_ (.A(_03011_),
    .B1(_12019_),
    .B2(_02748_),
    .ZN(_21813_));
 INV_X1 _38977_ (.A(_03155_),
    .ZN(_14127_));
 INV_X1 _38978_ (.A(_03147_),
    .ZN(_21839_));
 INV_X1 _38979_ (.A(_03154_),
    .ZN(_21843_));
 CLKBUF_X3 _38980_ (.A(_03272_),
    .Z(_12020_));
 AND2_X1 _38981_ (.A1(_00546_),
    .A2(_12020_),
    .ZN(_12021_));
 BUF_X4 _38982_ (.A(_03228_),
    .Z(_12022_));
 AOI21_X4 _38983_ (.A(_12021_),
    .B1(_12022_),
    .B2(_21883_),
    .ZN(_14134_));
 OAI21_X1 _38984_ (.A(_03557_),
    .B1(_03553_),
    .B2(_03560_),
    .ZN(_12023_));
 NAND2_X2 _38985_ (.A1(_03703_),
    .A2(_12023_),
    .ZN(_21957_));
 OR2_X1 _38986_ (.A1(_03533_),
    .A2(_21975_),
    .ZN(_12024_));
 AOI21_X1 _38987_ (.A(_03703_),
    .B1(_03842_),
    .B2(_12024_),
    .ZN(_12025_));
 AOI21_X1 _38988_ (.A(_12025_),
    .B1(_03703_),
    .B2(_21970_),
    .ZN(_21971_));
 CLKBUF_X3 _38989_ (.A(_03908_),
    .Z(_12026_));
 MUX2_X2 _38990_ (.A(_04197_),
    .B(_04199_),
    .S(_12026_),
    .Z(_14148_));
 AND2_X1 _38991_ (.A1(_00572_),
    .A2(_04566_),
    .ZN(_12027_));
 AOI21_X2 _38992_ (.A(_12027_),
    .B1(_12026_),
    .B2(_22006_),
    .ZN(_22044_));
 AND2_X1 _38993_ (.A1(_22003_),
    .A2(_12026_),
    .ZN(_12028_));
 AOI21_X2 _38994_ (.A(_12028_),
    .B1(_04566_),
    .B2(_00571_),
    .ZN(_22051_));
 AND2_X1 _38995_ (.A1(_22012_),
    .A2(_12026_),
    .ZN(_12029_));
 AOI21_X2 _38996_ (.A(_12029_),
    .B1(_04566_),
    .B2(_00569_),
    .ZN(_22058_));
 AND2_X1 _38997_ (.A1(_22015_),
    .A2(_12026_),
    .ZN(_12030_));
 AOI21_X2 _38998_ (.A(_12030_),
    .B1(_04566_),
    .B2(_00566_),
    .ZN(_22065_));
 AND2_X1 _38999_ (.A1(_22018_),
    .A2(_12026_),
    .ZN(_12031_));
 AOI21_X2 _39000_ (.A(_12031_),
    .B1(_04566_),
    .B2(_00567_),
    .ZN(_22072_));
 AND2_X1 _39001_ (.A1(_22021_),
    .A2(_12026_),
    .ZN(_12032_));
 AOI21_X2 _39002_ (.A(_12032_),
    .B1(_04566_),
    .B2(_00563_),
    .ZN(_22089_));
 INV_X1 _39003_ (.A(_04442_),
    .ZN(_22109_));
 CLKBUF_X3 _39004_ (.A(_04630_),
    .Z(_12033_));
 MUX2_X1 _39005_ (.A(_22168_),
    .B(_00574_),
    .S(_12033_),
    .Z(_12034_));
 INV_X2 _39006_ (.A(_12034_),
    .ZN(_14165_));
 MUX2_X1 _39007_ (.A(_22147_),
    .B(_00586_),
    .S(_12033_),
    .Z(_12035_));
 INV_X1 _39008_ (.A(_12035_),
    .ZN(_22191_));
 MUX2_X1 _39009_ (.A(_22153_),
    .B(_00583_),
    .S(_12033_),
    .Z(_12036_));
 INV_X1 _39010_ (.A(_12036_),
    .ZN(_22205_));
 MUX2_X1 _39011_ (.A(_22156_),
    .B(_00580_),
    .S(_12033_),
    .Z(_12037_));
 INV_X1 _39012_ (.A(_12037_),
    .ZN(_22212_));
 MUX2_X1 _39013_ (.A(_22165_),
    .B(_00578_),
    .S(_12033_),
    .Z(_12038_));
 INV_X1 _39014_ (.A(_12038_),
    .ZN(_22188_));
 MUX2_X1 _39015_ (.A(_22162_),
    .B(_00577_),
    .S(_12033_),
    .Z(_12039_));
 INV_X1 _39016_ (.A(_12039_),
    .ZN(_22236_));
 MUX2_X1 _39017_ (.A(_00575_),
    .B(_22171_),
    .S(_12033_),
    .Z(_12040_));
 INV_X1 _39018_ (.A(_12040_),
    .ZN(_22244_));
 BUF_X2 _39019_ (.A(_05406_),
    .Z(_12041_));
 AND2_X1 _39020_ (.A1(_00588_),
    .A2(_12041_),
    .ZN(_12042_));
 BUF_X4 _39021_ (.A(_05346_),
    .Z(_12043_));
 AOI21_X4 _39022_ (.A(_12042_),
    .B1(_12043_),
    .B2(_22315_),
    .ZN(_14182_));
 AND2_X1 _39023_ (.A1(_00600_),
    .A2(_12041_),
    .ZN(_12044_));
 AOI21_X2 _39024_ (.A(_12044_),
    .B1(_12043_),
    .B2(_22294_),
    .ZN(_22338_));
 AND2_X1 _39025_ (.A1(_00597_),
    .A2(_12041_),
    .ZN(_12045_));
 AOI21_X2 _39026_ (.A(_12045_),
    .B1(_12043_),
    .B2(_22300_),
    .ZN(_22352_));
 AND2_X1 _39027_ (.A1(_00594_),
    .A2(_12041_),
    .ZN(_12046_));
 AOI21_X2 _39028_ (.A(_12046_),
    .B1(_12043_),
    .B2(_22303_),
    .ZN(_22359_));
 AND2_X1 _39029_ (.A1(_00592_),
    .A2(_12041_),
    .ZN(_12047_));
 AOI21_X2 _39030_ (.A(_12047_),
    .B1(_12043_),
    .B2(_22312_),
    .ZN(_22335_));
 OAI21_X1 _39031_ (.A(_05685_),
    .B1(_05598_),
    .B2(_05597_),
    .ZN(_12048_));
 NOR2_X1 _39032_ (.A1(_05681_),
    .A2(_05609_),
    .ZN(_12049_));
 OAI21_X1 _39033_ (.A(_05853_),
    .B1(_05664_),
    .B2(_05621_),
    .ZN(_12050_));
 AOI21_X1 _39034_ (.A(_12048_),
    .B1(_12049_),
    .B2(_12050_),
    .ZN(_12051_));
 NAND2_X1 _39035_ (.A1(_05670_),
    .A2(_05593_),
    .ZN(_12052_));
 OAI21_X2 _39036_ (.A(_05716_),
    .B1(_12051_),
    .B2(_12052_),
    .ZN(_22395_));
 INV_X1 _39037_ (.A(_05937_),
    .ZN(_22409_));
 INV_X1 _39038_ (.A(_06034_),
    .ZN(_14189_));
 INV_X1 _39039_ (.A(_06022_),
    .ZN(_22421_));
 INV_X1 _39040_ (.A(_06033_),
    .ZN(_22425_));
 CLKBUF_X3 _39041_ (.A(_06102_),
    .Z(_12053_));
 MUX2_X1 _39042_ (.A(_22462_),
    .B(_00602_),
    .S(_12053_),
    .Z(_12054_));
 INV_X2 _39043_ (.A(_12054_),
    .ZN(_14196_));
 MUX2_X1 _39044_ (.A(_22441_),
    .B(_00614_),
    .S(_12053_),
    .Z(_12055_));
 INV_X1 _39045_ (.A(_12055_),
    .ZN(_22485_));
 MUX2_X1 _39046_ (.A(_22450_),
    .B(_00608_),
    .S(_12053_),
    .Z(_12056_));
 INV_X1 _39047_ (.A(_12056_),
    .ZN(_22506_));
 MUX2_X1 _39048_ (.A(_22459_),
    .B(_00606_),
    .S(_12053_),
    .Z(_12057_));
 INV_X1 _39049_ (.A(_12057_),
    .ZN(_22482_));
 MUX2_X1 _39050_ (.A(_22456_),
    .B(_00605_),
    .S(_12053_),
    .Z(_12058_));
 INV_X1 _39051_ (.A(_12058_),
    .ZN(_22530_));
 MUX2_X1 _39052_ (.A(_00603_),
    .B(_22465_),
    .S(_12053_),
    .Z(_12059_));
 INV_X1 _39053_ (.A(_12059_),
    .ZN(_22537_));
 OAI22_X2 _39054_ (.A1(_06478_),
    .A2(_06625_),
    .B1(_06651_),
    .B2(_06499_),
    .ZN(_22550_));
 INV_X1 _39055_ (.A(_22545_),
    .ZN(_22542_));
 XNOR2_X1 _39056_ (.A(_06547_),
    .B(_19424_),
    .ZN(_12060_));
 NOR2_X1 _39057_ (.A1(_06499_),
    .A2(_12060_),
    .ZN(_12061_));
 AOI21_X1 _39058_ (.A(_12061_),
    .B1(_06499_),
    .B2(_22555_),
    .ZN(_22557_));
 INV_X1 _39059_ (.A(_14205_),
    .ZN(_14210_));
 INV_X1 _39060_ (.A(_14225_),
    .ZN(_19482_));
 INV_X1 _39061_ (.A(_14224_),
    .ZN(_19487_));
 INV_X1 _39062_ (.A(_14244_),
    .ZN(_19539_));
 INV_X1 _39063_ (.A(_14243_),
    .ZN(_19544_));
 INV_X1 _39064_ (.A(_07049_),
    .ZN(_19552_));
 INV_X1 _39065_ (.A(_14263_),
    .ZN(_19596_));
 INV_X1 _39066_ (.A(_14262_),
    .ZN(_19601_));
 INV_X1 _39067_ (.A(_14276_),
    .ZN(_19653_));
 INV_X1 _39068_ (.A(_14294_),
    .ZN(_19710_));
 INV_X1 _39069_ (.A(_14311_),
    .ZN(_19767_));
 INV_X1 _39070_ (.A(_14333_),
    .ZN(_19824_));
 INV_X1 _39071_ (.A(_14332_),
    .ZN(_19829_));
 INV_X1 _39072_ (.A(_14350_),
    .ZN(_19881_));
 INV_X1 _39073_ (.A(_14362_),
    .ZN(_19938_));
 INV_X1 _39074_ (.A(_14384_),
    .ZN(_19995_));
 INV_X1 _39075_ (.A(_14383_),
    .ZN(_20000_));
 INV_X1 _39076_ (.A(_14396_),
    .ZN(_20052_));
 INV_X1 _39077_ (.A(_14418_),
    .ZN(_20109_));
 INV_X1 _39078_ (.A(_14417_),
    .ZN(_20114_));
 INV_X1 _39079_ (.A(_14430_),
    .ZN(_20166_));
 INV_X1 _39080_ (.A(_14434_),
    .ZN(_20171_));
 INV_X1 _39081_ (.A(_14447_),
    .ZN(_20223_));
 INV_X1 _39082_ (.A(_14469_),
    .ZN(_20280_));
 INV_X1 _39083_ (.A(_14468_),
    .ZN(_20285_));
 INV_X1 _39084_ (.A(_14486_),
    .ZN(_20337_));
 INV_X1 _39085_ (.A(_14485_),
    .ZN(_20342_));
 INV_X1 _39086_ (.A(_10424_),
    .ZN(_20395_));
 AND2_X1 _39087_ (.A1(_20362_),
    .A2(_11981_),
    .ZN(_12062_));
 AOI21_X2 _39088_ (.A(_12062_),
    .B1(_10394_),
    .B2(_00459_),
    .ZN(_20417_));
 AND2_X1 _39089_ (.A1(_20374_),
    .A2(_11981_),
    .ZN(_12063_));
 AOI21_X4 _39090_ (.A(_12063_),
    .B1(_10394_),
    .B2(_00454_),
    .ZN(_20431_));
 INV_X1 _39091_ (.A(_00456_),
    .ZN(_12064_));
 INV_X1 _39092_ (.A(_20368_),
    .ZN(_12065_));
 MUX2_X2 _39093_ (.A(_12064_),
    .B(_12065_),
    .S(_11981_),
    .Z(_20445_));
 AND2_X1 _39094_ (.A1(_20380_),
    .A2(_11981_),
    .ZN(_12066_));
 AOI21_X2 _39095_ (.A(_12066_),
    .B1(_10394_),
    .B2(_00451_),
    .ZN(_20455_));
 XNOR2_X1 _39096_ (.A(_10639_),
    .B(_20478_),
    .ZN(_12067_));
 NOR2_X1 _39097_ (.A1(_10795_),
    .A2(_12067_),
    .ZN(_12068_));
 AOI21_X1 _39098_ (.A(_12068_),
    .B1(_10795_),
    .B2(_20479_),
    .ZN(_20481_));
 AND2_X1 _39099_ (.A1(_11043_),
    .A2(_11045_),
    .ZN(_20539_));
 AND2_X1 _39100_ (.A1(_00462_),
    .A2(_11988_),
    .ZN(_12069_));
 AOI21_X4 _39101_ (.A(_12069_),
    .B1(_11991_),
    .B2(_20536_),
    .ZN(_14509_));
 AND2_X1 _39102_ (.A1(_00474_),
    .A2(_11988_),
    .ZN(_12070_));
 AOI21_X4 _39103_ (.A(_12070_),
    .B1(_11991_),
    .B2(_20515_),
    .ZN(_20554_));
 AND2_X1 _39104_ (.A1(_00473_),
    .A2(_11988_),
    .ZN(_12071_));
 AOI21_X4 _39105_ (.A(_12071_),
    .B1(_11991_),
    .B2(_20512_),
    .ZN(_20561_));
 NOR2_X1 _39106_ (.A1(_11097_),
    .A2(_11991_),
    .ZN(_12072_));
 AOI21_X2 _39107_ (.A(_12072_),
    .B1(_11991_),
    .B2(_20521_),
    .ZN(_20568_));
 NOR2_X1 _39108_ (.A1(_11108_),
    .A2(_11991_),
    .ZN(_12073_));
 AOI21_X2 _39109_ (.A(_12073_),
    .B1(_11991_),
    .B2(_20527_),
    .ZN(_20582_));
 XOR2_X1 _39110_ (.A(_11367_),
    .B(_20628_),
    .Z(_12074_));
 NAND2_X1 _39111_ (.A1(_11306_),
    .A2(_12074_),
    .ZN(_12075_));
 OAI21_X1 _39112_ (.A(_12075_),
    .B1(_11306_),
    .B2(_20623_),
    .ZN(_20625_));
 INV_X1 _39113_ (.A(_14578_),
    .ZN(_14574_));
 AND2_X1 _39114_ (.A1(_11722_),
    .A2(_11712_),
    .ZN(_20674_));
 INV_X1 _39115_ (.A(_14947_),
    .ZN(_14962_));
 AND2_X1 _39116_ (.A1(_11673_),
    .A2(_11754_),
    .ZN(_20708_));
 INV_X1 _39117_ (.A(_15164_),
    .ZN(_15161_));
 AND2_X1 _39118_ (.A1(_11698_),
    .A2(_11775_),
    .ZN(_20740_));
 AND2_X1 _39119_ (.A1(_11712_),
    .A2(_11774_),
    .ZN(_20751_));
 INV_X1 _39120_ (.A(_15654_),
    .ZN(_15656_));
 INV_X1 _39121_ (.A(_15967_),
    .ZN(_15977_));
 INV_X1 _39122_ (.A(_16463_),
    .ZN(_16490_));
 INV_X1 _39123_ (.A(_16516_),
    .ZN(_16499_));
 AND2_X1 _39124_ (.A1(_11698_),
    .A2(_11702_),
    .ZN(_20853_));
 INV_X1 _39125_ (.A(_17655_),
    .ZN(_18634_));
 INV_X1 _39126_ (.A(_16745_),
    .ZN(_16741_));
 INV_X1 _39127_ (.A(_16984_),
    .ZN(_16980_));
 INV_X1 _39128_ (.A(_18531_),
    .ZN(_17114_));
 INV_X1 _39129_ (.A(_17357_),
    .ZN(_17353_));
 INV_X1 _39130_ (.A(_17679_),
    .ZN(_17676_));
 INV_X1 _39131_ (.A(_18177_),
    .ZN(_18319_));
 INV_X1 _39132_ (.A(_18418_),
    .ZN(_18241_));
 MUX2_X1 _39133_ (.A(_00487_),
    .B(_21130_),
    .S(_11995_),
    .Z(_12076_));
 INV_X1 _39134_ (.A(_12076_),
    .ZN(_21179_));
 MUX2_X1 _39135_ (.A(_00485_),
    .B(_21139_),
    .S(_11995_),
    .Z(_12077_));
 INV_X1 _39136_ (.A(_12077_),
    .ZN(_21186_));
 MUX2_X1 _39137_ (.A(_00484_),
    .B(_21136_),
    .S(_11995_),
    .Z(_12078_));
 INV_X1 _39138_ (.A(_12078_),
    .ZN(_21207_));
 MUX2_X1 _39139_ (.A(_00480_),
    .B(_21151_),
    .S(_12193_),
    .Z(_12079_));
 INV_X1 _39140_ (.A(_12079_),
    .ZN(_21167_));
 MUX2_X1 _39141_ (.A(_12503_),
    .B(_12648_),
    .S(_12551_),
    .Z(_21237_));
 XNOR2_X1 _39142_ (.A(_12555_),
    .B(_21246_),
    .ZN(_12080_));
 NOR2_X1 _39143_ (.A1(_12644_),
    .A2(_12080_),
    .ZN(_12081_));
 AOI21_X1 _39144_ (.A(_12081_),
    .B1(_12644_),
    .B2(_21241_),
    .ZN(_21243_));
 INV_X1 _39145_ (.A(_12799_),
    .ZN(_21259_));
 NOR2_X1 _39146_ (.A1(_12937_),
    .A2(_12942_),
    .ZN(_21304_));
 MUX2_X2 _39147_ (.A(_12990_),
    .B(_12991_),
    .S(_13180_),
    .Z(_21319_));
 AND2_X1 _39148_ (.A1(_00501_),
    .A2(_12877_),
    .ZN(_12082_));
 AOI21_X2 _39149_ (.A(_12082_),
    .B1(_12004_),
    .B2(_21271_),
    .ZN(_21326_));
 NOR2_X1 _39150_ (.A1(_12963_),
    .A2(_12004_),
    .ZN(_12083_));
 AOI21_X4 _39151_ (.A(_12083_),
    .B1(_12004_),
    .B2(_21280_),
    .ZN(_21333_));
 AND2_X1 _39152_ (.A1(_00496_),
    .A2(_12877_),
    .ZN(_12084_));
 AOI21_X2 _39153_ (.A(_12084_),
    .B1(_12004_),
    .B2(_21283_),
    .ZN(_21340_));
 NOR2_X1 _39154_ (.A1(_12967_),
    .A2(_12004_),
    .ZN(_12085_));
 AOI21_X2 _39155_ (.A(_12085_),
    .B1(_12004_),
    .B2(_21286_),
    .ZN(_21347_));
 MUX2_X2 _39156_ (.A(_13022_),
    .B(_13023_),
    .S(_13180_),
    .Z(_21354_));
 NOR2_X1 _39157_ (.A1(_12978_),
    .A2(_12004_),
    .ZN(_12086_));
 AOI21_X2 _39158_ (.A(_12086_),
    .B1(_12004_),
    .B2(_21289_),
    .ZN(_21364_));
 NAND2_X2 _39159_ (.A1(_00683_),
    .A2(_00643_),
    .ZN(_21376_));
 AOI21_X1 _39160_ (.A(_00778_),
    .B1(_00779_),
    .B2(_00782_),
    .ZN(_21384_));
 XNOR2_X1 _39161_ (.A(_00658_),
    .B(_21387_),
    .ZN(_12087_));
 NOR2_X1 _39162_ (.A1(_00683_),
    .A2(_12087_),
    .ZN(_12088_));
 AOI21_X1 _39163_ (.A(_12088_),
    .B1(_00683_),
    .B2(_21388_),
    .ZN(_21390_));
 INV_X1 _39164_ (.A(_00910_),
    .ZN(_21402_));
 INV_X1 _39165_ (.A(_00917_),
    .ZN(_21406_));
 NOR3_X1 _39166_ (.A1(_00997_),
    .A2(_01069_),
    .A3(_12006_),
    .ZN(_12089_));
 NOR2_X1 _39167_ (.A1(_21448_),
    .A2(_01104_),
    .ZN(_12090_));
 AOI21_X1 _39168_ (.A(_12089_),
    .B1(_12090_),
    .B2(_00997_),
    .ZN(_21451_));
 MUX2_X1 _39169_ (.A(_01053_),
    .B(_01054_),
    .S(_12006_),
    .Z(_21466_));
 MUX2_X2 _39170_ (.A(_01056_),
    .B(_01057_),
    .S(_12006_),
    .Z(_21473_));
 AND2_X1 _39171_ (.A1(_21427_),
    .A2(_12006_),
    .ZN(_12091_));
 AOI21_X2 _39172_ (.A(_12091_),
    .B1(_01104_),
    .B2(_00513_),
    .ZN(_21480_));
 MUX2_X1 _39173_ (.A(_00510_),
    .B(_21430_),
    .S(_12006_),
    .Z(_12092_));
 INV_X1 _39174_ (.A(_12092_),
    .ZN(_21487_));
 AND2_X1 _39175_ (.A1(_21433_),
    .A2(_12006_),
    .ZN(_12093_));
 AOI21_X2 _39176_ (.A(_12093_),
    .B1(_01104_),
    .B2(_00511_),
    .ZN(_21494_));
 AND2_X1 _39177_ (.A1(_00512_),
    .A2(_01104_),
    .ZN(_12094_));
 AOI21_X2 _39178_ (.A(_12094_),
    .B1(_12006_),
    .B2(_21424_),
    .ZN(_21501_));
 MUX2_X1 _39179_ (.A(_00507_),
    .B(_21436_),
    .S(_00995_),
    .Z(_12095_));
 INV_X1 _39180_ (.A(_12095_),
    .ZN(_21511_));
 XNOR2_X1 _39181_ (.A(_01418_),
    .B(_21534_),
    .ZN(_12096_));
 NOR2_X1 _39182_ (.A1(_01597_),
    .A2(_12096_),
    .ZN(_12097_));
 AOI21_X1 _39183_ (.A(_12097_),
    .B1(_01597_),
    .B2(_21535_),
    .ZN(_21537_));
 MUX2_X1 _39184_ (.A(_00530_),
    .B(_21571_),
    .S(_12010_),
    .Z(_12098_));
 INV_X1 _39185_ (.A(_12098_),
    .ZN(_21610_));
 MUX2_X1 _39186_ (.A(_00529_),
    .B(_21568_),
    .S(_12010_),
    .Z(_12099_));
 INV_X1 _39187_ (.A(_12099_),
    .ZN(_21617_));
 MUX2_X1 _39188_ (.A(_00527_),
    .B(_21577_),
    .S(_12010_),
    .Z(_12100_));
 INV_X1 _39189_ (.A(_12100_),
    .ZN(_21624_));
 MUX2_X1 _39190_ (.A(_00524_),
    .B(_21580_),
    .S(_12010_),
    .Z(_12101_));
 INV_X1 _39191_ (.A(_12101_),
    .ZN(_21631_));
 MUX2_X1 _39192_ (.A(_00525_),
    .B(_21583_),
    .S(_12010_),
    .Z(_12102_));
 INV_X1 _39193_ (.A(_12102_),
    .ZN(_21638_));
 MUX2_X1 _39194_ (.A(_00526_),
    .B(_21574_),
    .S(_12010_),
    .Z(_12103_));
 INV_X1 _39195_ (.A(_12103_),
    .ZN(_21645_));
 MUX2_X1 _39196_ (.A(_00522_),
    .B(_21589_),
    .S(_01805_),
    .Z(_12104_));
 INV_X1 _39197_ (.A(_12104_),
    .ZN(_21606_));
 NOR2_X1 _39198_ (.A1(_02039_),
    .A2(_02092_),
    .ZN(_12105_));
 OAI21_X1 _39199_ (.A(_12105_),
    .B1(_02123_),
    .B2(_02150_),
    .ZN(_12106_));
 NAND2_X2 _39200_ (.A1(_02180_),
    .A2(_12106_),
    .ZN(_21667_));
 OAI21_X1 _39201_ (.A(_02224_),
    .B1(_02180_),
    .B2(_02261_),
    .ZN(_12107_));
 MUX2_X1 _39202_ (.A(_02085_),
    .B(_12107_),
    .S(_02196_),
    .Z(_21675_));
 NAND2_X1 _39203_ (.A1(_02174_),
    .A2(_21678_),
    .ZN(_12108_));
 NAND3_X1 _39204_ (.A1(_02207_),
    .A2(_02453_),
    .A3(_12108_),
    .ZN(_12109_));
 OAI21_X1 _39205_ (.A(_12109_),
    .B1(_02207_),
    .B2(_21679_),
    .ZN(_21681_));
 INV_X1 _39206_ (.A(_02452_),
    .ZN(_14113_));
 INV_X1 _39207_ (.A(_02444_),
    .ZN(_21693_));
 INV_X1 _39208_ (.A(_02451_),
    .ZN(_21697_));
 MUX2_X1 _39209_ (.A(_21712_),
    .B(_00544_),
    .S(_12014_),
    .Z(_12110_));
 INV_X1 _39210_ (.A(_12110_),
    .ZN(_21757_));
 MUX2_X1 _39211_ (.A(_21709_),
    .B(_00543_),
    .S(_12014_),
    .Z(_12111_));
 INV_X1 _39212_ (.A(_12111_),
    .ZN(_21764_));
 MUX2_X1 _39213_ (.A(_21718_),
    .B(_00541_),
    .S(_12014_),
    .Z(_12112_));
 INV_X1 _39214_ (.A(_12112_),
    .ZN(_21771_));
 MUX2_X1 _39215_ (.A(_21721_),
    .B(_00538_),
    .S(_12014_),
    .Z(_12113_));
 INV_X1 _39216_ (.A(_12113_),
    .ZN(_21778_));
 MUX2_X1 _39217_ (.A(_21724_),
    .B(_00539_),
    .S(_12014_),
    .Z(_12114_));
 INV_X1 _39218_ (.A(_12114_),
    .ZN(_21785_));
 MUX2_X1 _39219_ (.A(_21715_),
    .B(_00540_),
    .S(_12014_),
    .Z(_12115_));
 INV_X1 _39220_ (.A(_12115_),
    .ZN(_21792_));
 MUX2_X1 _39221_ (.A(_21727_),
    .B(_00535_),
    .S(_12014_),
    .Z(_12116_));
 INV_X1 _39222_ (.A(_12116_),
    .ZN(_21802_));
 XNOR2_X1 _39223_ (.A(_02920_),
    .B(_21825_),
    .ZN(_12117_));
 NOR2_X1 _39224_ (.A1(_03011_),
    .A2(_12117_),
    .ZN(_12118_));
 AOI21_X1 _39225_ (.A(_12118_),
    .B1(_03011_),
    .B2(_21826_),
    .ZN(_21828_));
 NOR3_X1 _39226_ (.A1(_03186_),
    .A2(_03259_),
    .A3(_12020_),
    .ZN(_12119_));
 AOI21_X1 _39227_ (.A(_12119_),
    .B1(_03260_),
    .B2(_12020_),
    .ZN(_21886_));
 AND2_X1 _39228_ (.A1(_00558_),
    .A2(_12020_),
    .ZN(_12120_));
 AOI21_X2 _39229_ (.A(_12120_),
    .B1(_12022_),
    .B2(_21862_),
    .ZN(_21901_));
 AND2_X1 _39230_ (.A1(_00557_),
    .A2(_12020_),
    .ZN(_12121_));
 AOI21_X2 _39231_ (.A(_12121_),
    .B1(_12022_),
    .B2(_21859_),
    .ZN(_21908_));
 AND2_X1 _39232_ (.A1(_21868_),
    .A2(_12022_),
    .ZN(_12122_));
 AOI21_X4 _39233_ (.A(_12122_),
    .B1(_12020_),
    .B2(_00555_),
    .ZN(_21915_));
 AND2_X1 _39234_ (.A1(_00552_),
    .A2(_12020_),
    .ZN(_12123_));
 AOI21_X4 _39235_ (.A(_12123_),
    .B1(_12022_),
    .B2(_21871_),
    .ZN(_21922_));
 MUX2_X1 _39236_ (.A(_00553_),
    .B(_21874_),
    .S(_12022_),
    .Z(_12124_));
 INV_X1 _39237_ (.A(_12124_),
    .ZN(_21929_));
 AND2_X1 _39238_ (.A1(_00554_),
    .A2(_12020_),
    .ZN(_12125_));
 AOI21_X2 _39239_ (.A(_12125_),
    .B1(_12022_),
    .B2(_21865_),
    .ZN(_21936_));
 AND2_X1 _39240_ (.A1(_00550_),
    .A2(_12020_),
    .ZN(_12126_));
 AOI21_X4 _39241_ (.A(_12126_),
    .B1(_12022_),
    .B2(_21880_),
    .ZN(_21897_));
 AND2_X1 _39242_ (.A1(_00549_),
    .A2(_12020_),
    .ZN(_12127_));
 AOI21_X2 _39243_ (.A(_12127_),
    .B1(_12022_),
    .B2(_21877_),
    .ZN(_21946_));
 AND2_X1 _39244_ (.A1(_00547_),
    .A2(_03272_),
    .ZN(_12128_));
 AOI21_X2 _39245_ (.A(_12128_),
    .B1(_12022_),
    .B2(_00548_),
    .ZN(_21953_));
 INV_X1 _39246_ (.A(_03841_),
    .ZN(_14144_));
 INV_X1 _39247_ (.A(_03833_),
    .ZN(_21984_));
 INV_X1 _39248_ (.A(_03840_),
    .ZN(_21988_));
 AOI21_X1 _39249_ (.A(_03963_),
    .B1(_03964_),
    .B2(_12026_),
    .ZN(_22030_));
 AND2_X1 _39250_ (.A1(_22009_),
    .A2(_12026_),
    .ZN(_12129_));
 AOI21_X2 _39251_ (.A(_12129_),
    .B1(_04566_),
    .B2(_00568_),
    .ZN(_22080_));
 MUX2_X2 _39252_ (.A(_04222_),
    .B(_04223_),
    .S(_12026_),
    .Z(_22041_));
 AND2_X1 _39253_ (.A1(_00562_),
    .A2(_03908_),
    .ZN(_12130_));
 AOI21_X2 _39254_ (.A(_12130_),
    .B1(_04566_),
    .B2(_00561_),
    .ZN(_22097_));
 NAND2_X1 _39255_ (.A1(_04182_),
    .A2(_04207_),
    .ZN(_12131_));
 AOI21_X1 _39256_ (.A(_04280_),
    .B1(_12131_),
    .B2(_04243_),
    .ZN(_12132_));
 NOR3_X1 _39257_ (.A1(_04156_),
    .A2(_04204_),
    .A3(_12132_),
    .ZN(_12133_));
 OAI21_X2 _39258_ (.A(_04312_),
    .B1(_12133_),
    .B2(_04239_),
    .ZN(_22102_));
 XNOR2_X1 _39259_ (.A(_04365_),
    .B(_22119_),
    .ZN(_12134_));
 NOR2_X1 _39260_ (.A1(_04312_),
    .A2(_12134_),
    .ZN(_12135_));
 AOI21_X1 _39261_ (.A(_12135_),
    .B1(_04312_),
    .B2(_22114_),
    .ZN(_22116_));
 INV_X1 _39262_ (.A(_14159_),
    .ZN(_14163_));
 INV_X1 _39263_ (.A(_04543_),
    .ZN(_22128_));
 INV_X1 _39264_ (.A(_04550_),
    .ZN(_22132_));
 MUX2_X1 _39265_ (.A(_22144_),
    .B(_00585_),
    .S(_12033_),
    .Z(_12136_));
 INV_X1 _39266_ (.A(_12136_),
    .ZN(_22199_));
 MUX2_X1 _39267_ (.A(_22159_),
    .B(_00581_),
    .S(_12033_),
    .Z(_12137_));
 INV_X1 _39268_ (.A(_12137_),
    .ZN(_22220_));
 MUX2_X1 _39269_ (.A(_22150_),
    .B(_00582_),
    .S(_12033_),
    .Z(_12138_));
 INV_X1 _39270_ (.A(_12138_),
    .ZN(_22227_));
 XNOR2_X1 _39271_ (.A(_05117_),
    .B(_22266_),
    .ZN(_12139_));
 NOR2_X1 _39272_ (.A1(_05084_),
    .A2(_12139_),
    .ZN(_12140_));
 AOI21_X1 _39273_ (.A(_12140_),
    .B1(_05084_),
    .B2(_22261_),
    .ZN(_22263_));
 AOI21_X1 _39274_ (.A(_05382_),
    .B1(_05378_),
    .B2(_12041_),
    .ZN(_22324_));
 AND2_X1 _39275_ (.A1(_00599_),
    .A2(_12041_),
    .ZN(_12141_));
 AOI21_X4 _39276_ (.A(_12141_),
    .B1(_12043_),
    .B2(_22291_),
    .ZN(_22346_));
 AND2_X1 _39277_ (.A1(_00595_),
    .A2(_12041_),
    .ZN(_12142_));
 AOI21_X2 _39278_ (.A(_12142_),
    .B1(_12043_),
    .B2(_22306_),
    .ZN(_22367_));
 AND2_X1 _39279_ (.A1(_00596_),
    .A2(_12041_),
    .ZN(_12143_));
 AOI21_X2 _39280_ (.A(_12143_),
    .B1(_12043_),
    .B2(_22297_),
    .ZN(_22374_));
 AND2_X1 _39281_ (.A1(_00591_),
    .A2(_12041_),
    .ZN(_12144_));
 AOI21_X2 _39282_ (.A(_12144_),
    .B1(_12043_),
    .B2(_22309_),
    .ZN(_22384_));
 AND2_X1 _39283_ (.A1(_22318_),
    .A2(_05406_),
    .ZN(_12145_));
 AOI21_X2 _39284_ (.A(_12145_),
    .B1(_12043_),
    .B2(_00589_),
    .ZN(_22391_));
 INV_X1 _39285_ (.A(_05911_),
    .ZN(_22404_));
 XNOR2_X1 _39286_ (.A(_05714_),
    .B(_22407_),
    .ZN(_12146_));
 NAND2_X1 _39287_ (.A1(_05746_),
    .A2(_12146_),
    .ZN(_12147_));
 OAI21_X1 _39288_ (.A(_12147_),
    .B1(_05746_),
    .B2(_22408_),
    .ZN(_22410_));
 MUX2_X1 _39289_ (.A(_22438_),
    .B(_00613_),
    .S(_12053_),
    .Z(_12148_));
 INV_X1 _39290_ (.A(_12148_),
    .ZN(_22493_));
 MUX2_X1 _39291_ (.A(_22447_),
    .B(_00611_),
    .S(_12053_),
    .Z(_12149_));
 INV_X1 _39292_ (.A(_12149_),
    .ZN(_22500_));
 MUX2_X1 _39293_ (.A(_22453_),
    .B(_00609_),
    .S(_12053_),
    .Z(_12150_));
 INV_X1 _39294_ (.A(_12150_),
    .ZN(_22514_));
 MUX2_X1 _39295_ (.A(_22444_),
    .B(_00610_),
    .S(_12053_),
    .Z(_12151_));
 INV_X1 _39296_ (.A(_12151_),
    .ZN(_22521_));
 NAND2_X2 _39297_ (.A1(_06499_),
    .A2(_06474_),
    .ZN(_22543_));
 INV_X1 _39298_ (.A(_20675_),
    .ZN(_14696_));
 INV_X1 _39299_ (.A(_20710_),
    .ZN(_15019_));
 INV_X1 _39300_ (.A(_20742_),
    .ZN(_15382_));
 INV_X1 _39301_ (.A(_20753_),
    .ZN(_15459_));
 INV_X1 _39302_ (.A(_20764_),
    .ZN(_15603_));
 INV_X1 _39303_ (.A(_20802_),
    .ZN(_16130_));
 INV_X1 _39304_ (.A(_20855_),
    .ZN(_16548_));
 INV_X1 _39305_ (.A(_20873_),
    .ZN(_17936_));
 INV_X1 _39306_ (.A(_20881_),
    .ZN(_16653_));
 INV_X1 _39307_ (.A(_19486_),
    .ZN(_14227_));
 INV_X1 _39308_ (.A(_19543_),
    .ZN(_14246_));
 INV_X1 _39309_ (.A(_19600_),
    .ZN(_14264_));
 INV_X1 _39310_ (.A(_19657_),
    .ZN(_14284_));
 INV_X1 _39311_ (.A(_19714_),
    .ZN(_14300_));
 INV_X1 _39312_ (.A(_19771_),
    .ZN(_14317_));
 INV_X1 _39313_ (.A(_19828_),
    .ZN(_14335_));
 INV_X1 _39314_ (.A(_19885_),
    .ZN(_14352_));
 INV_X1 _39315_ (.A(_19942_),
    .ZN(_14369_));
 INV_X1 _39316_ (.A(_19999_),
    .ZN(_14385_));
 INV_X1 _39317_ (.A(_20056_),
    .ZN(_14402_));
 INV_X1 _39318_ (.A(_20113_),
    .ZN(_14419_));
 INV_X1 _39319_ (.A(_20170_),
    .ZN(_14436_));
 INV_X1 _39320_ (.A(_20227_),
    .ZN(_14454_));
 INV_X1 _39321_ (.A(_20284_),
    .ZN(_14471_));
 INV_X1 _39322_ (.A(_20341_),
    .ZN(_14487_));
 INV_X1 _39323_ (.A(_20646_),
    .ZN(_14523_));
 INV_X1 _39324_ (.A(_20651_),
    .ZN(_14586_));
 INV_X1 _39325_ (.A(_20656_),
    .ZN(_14616_));
 INV_X1 _39326_ (.A(_19087_),
    .ZN(_19083_));
 INV_X1 _39327_ (.A(_20665_),
    .ZN(_19077_));
 INV_X1 _39328_ (.A(_20668_),
    .ZN(_19402_));
 INV_X1 _39329_ (.A(_20671_),
    .ZN(_14652_));
 INV_X1 _39330_ (.A(_19412_),
    .ZN(_19408_));
 INV_X1 _39331_ (.A(_20685_),
    .ZN(_14721_));
 INV_X1 _39332_ (.A(_20691_),
    .ZN(_14760_));
 INV_X1 _39333_ (.A(_20694_),
    .ZN(_14780_));
 INV_X1 _39334_ (.A(_20706_),
    .ZN(_15683_));
 INV_X1 _39335_ (.A(_20713_),
    .ZN(_15673_));
 INV_X1 _39336_ (.A(_20717_),
    .ZN(_15059_));
 INV_X1 _39337_ (.A(_20723_),
    .ZN(_15311_));
 INV_X1 _39338_ (.A(_20726_),
    .ZN(_19213_));
 INV_X1 _39339_ (.A(_20729_),
    .ZN(_19359_));
 INV_X1 _39340_ (.A(_20735_),
    .ZN(_19364_));
 INV_X1 _39341_ (.A(_20746_),
    .ZN(_15401_));
 INV_X1 _39342_ (.A(_20749_),
    .ZN(_15448_));
 INV_X1 _39343_ (.A(_20756_),
    .ZN(_19220_));
 INV_X1 _39344_ (.A(_20759_),
    .ZN(_15505_));
 INV_X1 _39345_ (.A(_20769_),
    .ZN(_19308_));
 INV_X1 _39346_ (.A(_19318_),
    .ZN(_19314_));
 INV_X1 _39347_ (.A(_20777_),
    .ZN(_15732_));
 INV_X1 _39348_ (.A(_20783_),
    .ZN(_15792_));
 INV_X1 _39349_ (.A(_20786_),
    .ZN(_15806_));
 INV_X1 _39350_ (.A(_20792_),
    .ZN(_15866_));
 INV_X1 _39351_ (.A(_20798_),
    .ZN(_16101_));
 INV_X1 _39352_ (.A(_20806_),
    .ZN(_16180_));
 INV_X1 _39353_ (.A(_20811_),
    .ZN(_16207_));
 INV_X1 _39354_ (.A(_20815_),
    .ZN(_19131_));
 INV_X1 _39355_ (.A(_20822_),
    .ZN(_19258_));
 INV_X1 _39356_ (.A(_19268_),
    .ZN(_19264_));
 INV_X1 _39357_ (.A(_20830_),
    .ZN(_16241_));
 INV_X1 _39358_ (.A(_20837_),
    .ZN(_16280_));
 INV_X1 _39359_ (.A(_20840_),
    .ZN(_19171_));
 INV_X1 _39360_ (.A(_20843_),
    .ZN(_16294_));
 INV_X1 _39361_ (.A(_20849_),
    .ZN(_16358_));
 INV_X1 _39362_ (.A(_20859_),
    .ZN(_16535_));
 INV_X1 _39363_ (.A(_20863_),
    .ZN(_19177_));
 INV_X1 _39364_ (.A(_20869_),
    .ZN(_16628_));
 INV_X1 _39365_ (.A(_20878_),
    .ZN(_18601_));
 INV_X1 _39366_ (.A(_20887_),
    .ZN(_18722_));
 INV_X1 _39367_ (.A(_20890_),
    .ZN(_16734_));
 INV_X1 _39368_ (.A(_20895_),
    .ZN(_17514_));
 INV_X1 _39369_ (.A(_20900_),
    .ZN(_18446_));
 INV_X1 _39370_ (.A(_20904_),
    .ZN(_16843_));
 INV_X1 _39371_ (.A(_20907_),
    .ZN(_18436_));
 INV_X1 _39372_ (.A(_20913_),
    .ZN(_16904_));
 INV_X1 _39373_ (.A(_20920_),
    .ZN(_17566_));
 INV_X1 _39374_ (.A(_20923_),
    .ZN(_16968_));
 INV_X1 _39375_ (.A(_20930_),
    .ZN(_17064_));
 INV_X1 _39376_ (.A(_20934_),
    .ZN(_18549_));
 INV_X1 _39377_ (.A(_18863_),
    .ZN(_18860_));
 INV_X1 _39378_ (.A(_20942_),
    .ZN(_17189_));
 INV_X1 _39379_ (.A(_20948_),
    .ZN(_17202_));
 INV_X1 _39380_ (.A(_20953_),
    .ZN(_18499_));
 INV_X1 _39381_ (.A(_18818_),
    .ZN(_18814_));
 INV_X1 _39382_ (.A(_20962_),
    .ZN(_18658_));
 INV_X1 _39383_ (.A(_20966_),
    .ZN(_17275_));
 INV_X1 _39384_ (.A(_20971_),
    .ZN(_17307_));
 INV_X1 _39385_ (.A(_20978_),
    .ZN(_18651_));
 INV_X1 _39386_ (.A(_20985_),
    .ZN(_19038_));
 INV_X1 _39387_ (.A(_20990_),
    .ZN(_17501_));
 INV_X1 _39388_ (.A(_20994_),
    .ZN(_17866_));
 INV_X1 _39389_ (.A(_20997_),
    .ZN(_17543_));
 INV_X1 _39390_ (.A(_21003_),
    .ZN(_18767_));
 INV_X1 _39391_ (.A(_21011_),
    .ZN(_17788_));
 INV_X1 _39392_ (.A(_21017_),
    .ZN(_18328_));
 INV_X1 _39393_ (.A(_21024_),
    .ZN(_17916_));
 INV_X1 _39394_ (.A(_21027_),
    .ZN(_18286_));
 INV_X1 _39395_ (.A(_21031_),
    .ZN(_18166_));
 INV_X1 _39396_ (.A(_21036_),
    .ZN(_18492_));
 INV_X1 _39397_ (.A(_21040_),
    .ZN(_18541_));
 INV_X1 _39398_ (.A(_21046_),
    .ZN(_18116_));
 INV_X1 _39399_ (.A(_21050_),
    .ZN(_18954_));
 INV_X1 _39400_ (.A(_21053_),
    .ZN(_18335_));
 INV_X1 _39401_ (.A(_21056_),
    .ZN(_18593_));
 INV_X1 _39402_ (.A(_21067_),
    .ZN(_18996_));
 INV_X1 _39403_ (.A(_21074_),
    .ZN(_18908_));
 INV_X1 _39404_ (.A(_20647_),
    .ZN(_14541_));
 INV_X1 _39405_ (.A(_20672_),
    .ZN(_14653_));
 INV_X1 _39406_ (.A(_20702_),
    .ZN(_15310_));
 INV_X1 _39407_ (.A(_20709_),
    .ZN(_15058_));
 INV_X1 _39408_ (.A(_20741_),
    .ZN(_15400_));
 INV_X1 _39409_ (.A(_20752_),
    .ZN(_15504_));
 INV_X1 _39410_ (.A(_20714_),
    .ZN(_15674_));
 INV_X1 _39411_ (.A(_20789_),
    .ZN(_15865_));
 INV_X1 _39412_ (.A(_20799_),
    .ZN(_16100_));
 INV_X1 _39413_ (.A(_20836_),
    .ZN(_16313_));
 INV_X1 _39414_ (.A(_20846_),
    .ZN(_16357_));
 INV_X1 _39415_ (.A(_20854_),
    .ZN(_16533_));
 INV_X1 _39416_ (.A(_20870_),
    .ZN(_16627_));
 INV_X1 _39417_ (.A(_20874_),
    .ZN(_17935_));
 INV_X1 _39418_ (.A(_20901_),
    .ZN(_18447_));
 INV_X1 _39419_ (.A(_20916_),
    .ZN(_18115_));
 INV_X1 _39420_ (.A(_20943_),
    .ZN(_17188_));
 INV_X1 _39421_ (.A(_20949_),
    .ZN(_17214_));
 INV_X1 _39422_ (.A(_20965_),
    .ZN(_17308_));
 INV_X1 _39423_ (.A(_20991_),
    .ZN(_17500_));
 INV_X1 _39424_ (.A(_20896_),
    .ZN(_17515_));
 INV_X1 _39425_ (.A(_21028_),
    .ZN(_18287_));
 AND2_X1 _39426_ (.A1(_11857_),
    .A2(_11685_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39427_ (.A1(_11665_),
    .A2(_11685_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39428_ (.A1(_11857_),
    .A2(_11884_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t1[2] ));
 BUF_X1 _39429_ (.A(_11667_),
    .Z(_12152_));
 AND2_X1 _39430_ (.A1(_12152_),
    .A2(_11686_),
    .ZN(\g_row[0].g_col[0].mult.stage1.dadda.t2[1] ));
 BUF_X1 _39431_ (.A(_11803_),
    .Z(_12153_));
 AND2_X1 _39432_ (.A1(_11764_),
    .A2(_12153_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39433_ (.A1(_11764_),
    .A2(_11765_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39434_ (.A1(_11851_),
    .A2(_11948_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39435_ (.A1(_11767_),
    .A2(_12153_),
    .ZN(\g_row[0].g_col[1].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39436_ (.A1(_11946_),
    .A2(_11771_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39437_ (.A1(_11873_),
    .A2(_11771_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39438_ (.A1(_11946_),
    .A2(_11940_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39439_ (.A1(_11946_),
    .A2(_11773_),
    .ZN(\g_row[0].g_col[2].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39440_ (.A1(_11781_),
    .A2(_11795_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39441_ (.A1(_11931_),
    .A2(_11795_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39442_ (.A1(_11781_),
    .A2(_11924_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39443_ (.A1(_11781_),
    .A2(_11794_),
    .ZN(\g_row[0].g_col[3].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39444_ (.A1(_12152_),
    .A2(_11814_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39445_ (.A1(_11665_),
    .A2(_11814_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39446_ (.A1(_12152_),
    .A2(_11915_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39447_ (.A1(_12152_),
    .A2(_11813_),
    .ZN(\g_row[1].g_col[0].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39448_ (.A1(_11851_),
    .A2(_11847_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39449_ (.A1(_11765_),
    .A2(_11847_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39450_ (.A1(_12153_),
    .A2(_11903_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39451_ (.A1(_12153_),
    .A2(_11846_),
    .ZN(\g_row[1].g_col[1].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39452_ (.A1(_11946_),
    .A2(_11872_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39453_ (.A1(_11873_),
    .A2(_11872_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39454_ (.A1(_11875_),
    .A2(_11958_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39455_ (.A1(_11875_),
    .A2(_11871_),
    .ZN(\g_row[1].g_col[2].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39456_ (.A1(_11761_),
    .A2(_11876_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39457_ (.A1(_11931_),
    .A2(_11876_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39458_ (.A1(_11761_),
    .A2(_11960_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39459_ (.A1(_11761_),
    .A2(_11877_),
    .ZN(\g_row[1].g_col[3].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39460_ (.A1(_11642_),
    .A2(_12152_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39461_ (.A1(_11665_),
    .A2(_11642_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39462_ (.A1(_12152_),
    .A2(_11649_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39463_ (.A1(_11644_),
    .A2(_12152_),
    .ZN(\g_row[2].g_col[0].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39464_ (.A1(_12153_),
    .A2(_11844_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39465_ (.A1(_11765_),
    .A2(_11844_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39466_ (.A1(_12153_),
    .A2(_11840_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39467_ (.A1(_12153_),
    .A2(_11843_),
    .ZN(\g_row[2].g_col[1].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39468_ (.A1(_11722_),
    .A2(_11875_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39469_ (.A1(_11722_),
    .A2(_11718_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39470_ (.A1(_11711_),
    .A2(_11875_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39471_ (.A1(_11702_),
    .A2(_11875_),
    .ZN(\g_row[2].g_col[2].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39472_ (.A1(_11761_),
    .A2(_11754_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39473_ (.A1(_11931_),
    .A2(_11754_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39474_ (.A1(_11761_),
    .A2(_11753_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39475_ (.A1(_11761_),
    .A2(_11755_),
    .ZN(\g_row[2].g_col[3].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39476_ (.A1(_12152_),
    .A2(_11854_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39477_ (.A1(_11665_),
    .A2(_11854_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39478_ (.A1(_12152_),
    .A2(_11856_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39479_ (.A1(_12152_),
    .A2(_11855_),
    .ZN(\g_row[3].g_col[0].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39480_ (.A1(_11799_),
    .A2(_12153_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39481_ (.A1(_11765_),
    .A2(_11799_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39482_ (.A1(_11806_),
    .A2(_12153_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39483_ (.A1(_11798_),
    .A2(_12153_),
    .ZN(\g_row[3].g_col[1].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39484_ (.A1(_11875_),
    .A2(_11774_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39485_ (.A1(_11873_),
    .A2(_11774_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39486_ (.A1(_11875_),
    .A2(_11779_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39487_ (.A1(_11875_),
    .A2(_11775_),
    .ZN(\g_row[3].g_col[2].mult.stage1.dadda.t2[1] ));
 AND2_X1 _39488_ (.A1(_11689_),
    .A2(_11761_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[0] ));
 AND2_X1 _39489_ (.A1(_11931_),
    .A2(_11689_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[1] ));
 AND2_X1 _39490_ (.A1(_11731_),
    .A2(_11761_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t1[2] ));
 AND2_X1 _39491_ (.A1(_11687_),
    .A2(_11761_),
    .ZN(\g_row[3].g_col[3].mult.stage1.dadda.t2[1] ));
 FA_X1 _39492_ (.A(_14058_),
    .B(_14059_),
    .CI(_14060_),
    .CO(_14061_),
    .S(_14062_));
 FA_X1 _39493_ (.A(_14060_),
    .B(_14063_),
    .CI(_14064_),
    .CO(_14065_),
    .S(_14066_));
 FA_X1 _39494_ (.A(_14067_),
    .B(_14068_),
    .CI(_14069_),
    .CO(_14070_),
    .S(_14071_));
 FA_X1 _39495_ (.A(_14073_),
    .B(_14074_),
    .CI(_14075_),
    .CO(_14076_),
    .S(_14077_));
 FA_X1 _39496_ (.A(_14075_),
    .B(_14078_),
    .CI(_14079_),
    .CO(_14080_),
    .S(_14081_));
 FA_X1 _39497_ (.A(_14082_),
    .B(_14083_),
    .CI(_14084_),
    .CO(_14085_),
    .S(_14086_));
 FA_X1 _39498_ (.A(_14088_),
    .B(_14089_),
    .CI(_14090_),
    .CO(_14091_),
    .S(_14092_));
 FA_X1 _39499_ (.A(_14090_),
    .B(_14093_),
    .CI(_14094_),
    .CO(_14095_),
    .S(_14096_));
 FA_X1 _39500_ (.A(_14097_),
    .B(_14098_),
    .CI(_14099_),
    .CO(_14100_),
    .S(_14101_));
 FA_X1 _39501_ (.A(_14103_),
    .B(_14104_),
    .CI(_14105_),
    .CO(_14106_),
    .S(_14107_));
 FA_X1 _39502_ (.A(_14105_),
    .B(_14108_),
    .CI(_14109_),
    .CO(_14110_),
    .S(_14111_));
 FA_X1 _39503_ (.A(_14112_),
    .B(_14113_),
    .CI(_14114_),
    .CO(_14115_),
    .S(_14116_));
 FA_X1 _39504_ (.A(_14118_),
    .B(_14119_),
    .CI(_14120_),
    .CO(_14121_),
    .S(_14122_));
 FA_X1 _39505_ (.A(_14120_),
    .B(_14123_),
    .CI(_14124_),
    .CO(_14125_),
    .S(_14126_));
 FA_X1 _39506_ (.A(_14127_),
    .B(_14128_),
    .CI(_14129_),
    .CO(_14130_),
    .S(_14131_));
 FA_X1 _39507_ (.A(_14133_),
    .B(_14134_),
    .CI(_14135_),
    .CO(_14136_),
    .S(_14137_));
 FA_X1 _39508_ (.A(_14134_),
    .B(_14138_),
    .CI(_14139_),
    .CO(_14140_),
    .S(_14141_));
 FA_X1 _39509_ (.A(_14142_),
    .B(_14143_),
    .CI(_14144_),
    .CO(_14145_),
    .S(_14146_));
 FA_X1 _39510_ (.A(_14148_),
    .B(_14149_),
    .CI(_14150_),
    .CO(_14151_),
    .S(_14152_));
 FA_X1 _39511_ (.A(_14148_),
    .B(_14153_),
    .CI(_14154_),
    .CO(_14155_),
    .S(_14156_));
 FA_X1 _39512_ (.A(_14157_),
    .B(_14158_),
    .CI(_14159_),
    .CO(_14160_),
    .S(_14161_));
 FA_X1 _39513_ (.A(_14164_),
    .B(_14165_),
    .CI(_14166_),
    .CO(_14167_),
    .S(_14168_));
 FA_X1 _39514_ (.A(_14165_),
    .B(_14169_),
    .CI(_14170_),
    .CO(_14171_),
    .S(_14172_));
 FA_X1 _39515_ (.A(_14173_),
    .B(_14174_),
    .CI(_14175_),
    .CO(_14176_),
    .S(_14177_));
 FA_X1 _39516_ (.A(_14180_),
    .B(_14181_),
    .CI(_14182_),
    .CO(_14183_),
    .S(_14184_));
 FA_X1 _39517_ (.A(_14182_),
    .B(_14185_),
    .CI(_14186_),
    .CO(_14187_),
    .S(_14188_));
 FA_X1 _39518_ (.A(_14189_),
    .B(_14190_),
    .CI(_14191_),
    .CO(_14192_),
    .S(_14193_));
 FA_X1 _39519_ (.A(_14195_),
    .B(_14196_),
    .CI(_14197_),
    .CO(_14198_),
    .S(_14199_));
 FA_X1 _39520_ (.A(_14196_),
    .B(_14200_),
    .CI(_14201_),
    .CO(_14202_),
    .S(_14203_));
 FA_X1 _39521_ (.A(_14204_),
    .B(_14205_),
    .CI(_14206_),
    .CO(_14207_),
    .S(_14208_));
 FA_X1 _39522_ (.A(_14211_),
    .B(_14212_),
    .CI(_14213_),
    .CO(_14214_),
    .S(_14215_));
 FA_X1 _39523_ (.A(_14216_),
    .B(_14217_),
    .CI(_14218_),
    .CO(_14219_),
    .S(_14220_));
 FA_X1 _39524_ (.A(_14222_),
    .B(_14223_),
    .CI(_14221_),
    .CO(_14224_),
    .S(_14225_));
 FA_X1 _39525_ (.A(_14226_),
    .B(_14227_),
    .CI(_14224_),
    .CO(_14228_),
    .S(_14229_));
 FA_X1 _39526_ (.A(_14230_),
    .B(_14231_),
    .CI(_14232_),
    .CO(_14233_),
    .S(_14234_));
 FA_X1 _39527_ (.A(_14235_),
    .B(_14236_),
    .CI(_14237_),
    .CO(_14238_),
    .S(_14239_));
 FA_X1 _39528_ (.A(_14241_),
    .B(_14242_),
    .CI(_14240_),
    .CO(_14243_),
    .S(_14244_));
 FA_X1 _39529_ (.A(_14245_),
    .B(_14246_),
    .CI(_14243_),
    .CO(_14247_),
    .S(_14248_));
 FA_X1 _39530_ (.A(_14249_),
    .B(_14250_),
    .CI(_14251_),
    .CO(_14252_),
    .S(_14253_));
 FA_X1 _39531_ (.A(_14254_),
    .B(_14255_),
    .CI(_14256_),
    .CO(_14257_),
    .S(_14258_));
 FA_X1 _39532_ (.A(_14259_),
    .B(_14260_),
    .CI(_14261_),
    .CO(_14262_),
    .S(_14263_));
 FA_X1 _39533_ (.A(_14264_),
    .B(_14262_),
    .CI(_14265_),
    .CO(_14266_),
    .S(_14267_));
 FA_X1 _39534_ (.A(_14268_),
    .B(_14269_),
    .CI(_14270_),
    .CO(_14271_),
    .S(_14272_));
 FA_X1 _39535_ (.A(_14273_),
    .B(_14274_),
    .CI(_14275_),
    .CO(_14276_),
    .S(_14277_));
 FA_X1 _39536_ (.A(_14278_),
    .B(_14279_),
    .CI(_14280_),
    .CO(_14281_),
    .S(_14282_));
 FA_X1 _39537_ (.A(_14283_),
    .B(_14281_),
    .CI(_14284_),
    .CO(_14285_),
    .S(_14286_));
 FA_X1 _39538_ (.A(_14287_),
    .B(_14288_),
    .CI(_14289_),
    .CO(_14290_),
    .S(_14291_));
 FA_X1 _39539_ (.A(_14216_),
    .B(_14292_),
    .CI(_14293_),
    .CO(_14294_),
    .S(_14295_));
 FA_X1 _39540_ (.A(_14222_),
    .B(_14296_),
    .CI(_14297_),
    .CO(_14298_),
    .S(_14299_));
 FA_X1 _39541_ (.A(_14298_),
    .B(_14300_),
    .CI(_14301_),
    .CO(_14302_),
    .S(_14303_));
 FA_X1 _39542_ (.A(_14304_),
    .B(_14305_),
    .CI(_14306_),
    .CO(_14307_),
    .S(_14308_));
 FA_X1 _39543_ (.A(_14235_),
    .B(_14309_),
    .CI(_14310_),
    .CO(_14311_),
    .S(_14312_));
 FA_X1 _39544_ (.A(_14241_),
    .B(_14313_),
    .CI(_14314_),
    .CO(_14315_),
    .S(_14316_));
 FA_X1 _39545_ (.A(_14315_),
    .B(_14317_),
    .CI(_14318_),
    .CO(_14319_),
    .S(_14320_));
 FA_X1 _39546_ (.A(_14321_),
    .B(_14322_),
    .CI(_14323_),
    .CO(_14324_),
    .S(_14325_));
 FA_X1 _39547_ (.A(_14254_),
    .B(_14326_),
    .CI(_14327_),
    .CO(_14328_),
    .S(_14329_));
 FA_X1 _39548_ (.A(_14259_),
    .B(_14331_),
    .CI(_14330_),
    .CO(_14332_),
    .S(_14333_));
 FA_X1 _39549_ (.A(_14334_),
    .B(_14335_),
    .CI(_14332_),
    .CO(_14336_),
    .S(_14337_));
 FA_X1 _39550_ (.A(_14338_),
    .B(_14339_),
    .CI(_14340_),
    .CO(_14341_),
    .S(_14342_));
 FA_X1 _39551_ (.A(_14273_),
    .B(_14343_),
    .CI(_14344_),
    .CO(_14345_),
    .S(_14346_));
 FA_X1 _39552_ (.A(_14278_),
    .B(_14348_),
    .CI(_14347_),
    .CO(_14349_),
    .S(_14350_));
 FA_X1 _39553_ (.A(_14349_),
    .B(_14351_),
    .CI(_14352_),
    .CO(_14353_),
    .S(_14354_));
 FA_X1 _39554_ (.A(_14355_),
    .B(_14356_),
    .CI(_14357_),
    .CO(_14358_),
    .S(_14359_));
 FA_X1 _39555_ (.A(_14216_),
    .B(_14360_),
    .CI(_14361_),
    .CO(_14362_),
    .S(_14363_));
 FA_X1 _39556_ (.A(_14222_),
    .B(_14364_),
    .CI(_14365_),
    .CO(_14366_),
    .S(_14367_));
 FA_X1 _39557_ (.A(_14368_),
    .B(_14366_),
    .CI(_14369_),
    .CO(_14370_),
    .S(_14371_));
 FA_X1 _39558_ (.A(_14372_),
    .B(_14373_),
    .CI(_14374_),
    .CO(_14375_),
    .S(_14376_));
 FA_X1 _39559_ (.A(_14235_),
    .B(_14377_),
    .CI(_14378_),
    .CO(_14379_),
    .S(_14380_));
 FA_X1 _39560_ (.A(_14241_),
    .B(_14381_),
    .CI(_14382_),
    .CO(_14383_),
    .S(_14384_));
 FA_X1 _39561_ (.A(_14385_),
    .B(_14383_),
    .CI(_14386_),
    .CO(_14387_),
    .S(_14388_));
 FA_X1 _39562_ (.A(_14389_),
    .B(_14390_),
    .CI(_14391_),
    .CO(_14392_),
    .S(_14393_));
 FA_X1 _39563_ (.A(_14254_),
    .B(_14394_),
    .CI(_14395_),
    .CO(_14396_),
    .S(_14397_));
 FA_X1 _39564_ (.A(_14259_),
    .B(_14399_),
    .CI(_14398_),
    .CO(_14400_),
    .S(_14401_));
 FA_X1 _39565_ (.A(_14400_),
    .B(_14402_),
    .CI(_14403_),
    .CO(_14404_),
    .S(_14405_));
 FA_X1 _39566_ (.A(_14406_),
    .B(_14407_),
    .CI(_14408_),
    .CO(_14409_),
    .S(_14410_));
 FA_X1 _39567_ (.A(_14273_),
    .B(_14411_),
    .CI(_14412_),
    .CO(_14413_),
    .S(_14414_));
 FA_X1 _39568_ (.A(_14278_),
    .B(_14415_),
    .CI(_14416_),
    .CO(_14417_),
    .S(_14418_));
 FA_X1 _39569_ (.A(_14419_),
    .B(_14417_),
    .CI(_14420_),
    .CO(_14421_),
    .S(_14422_));
 FA_X1 _39570_ (.A(_14423_),
    .B(_14424_),
    .CI(_14425_),
    .CO(_14426_),
    .S(_14427_));
 FA_X1 _39571_ (.A(_14216_),
    .B(_14428_),
    .CI(_14429_),
    .CO(_14430_),
    .S(_14431_));
 FA_X1 _39572_ (.A(_14222_),
    .B(_14432_),
    .CI(_14433_),
    .CO(_14434_),
    .S(_14435_));
 FA_X1 _39573_ (.A(_14436_),
    .B(_14434_),
    .CI(_14437_),
    .CO(_14438_),
    .S(_14439_));
 FA_X1 _39574_ (.A(_14440_),
    .B(_14441_),
    .CI(_14442_),
    .CO(_14443_),
    .S(_14444_));
 FA_X1 _39575_ (.A(_14235_),
    .B(_14445_),
    .CI(_14446_),
    .CO(_14447_),
    .S(_14448_));
 FA_X1 _39576_ (.A(_14241_),
    .B(_14449_),
    .CI(_14450_),
    .CO(_14451_),
    .S(_14452_));
 FA_X1 _39577_ (.A(_14453_),
    .B(_14451_),
    .CI(_14454_),
    .CO(_14455_),
    .S(_14456_));
 FA_X1 _39578_ (.A(_14457_),
    .B(_14458_),
    .CI(_14459_),
    .CO(_14460_),
    .S(_14461_));
 FA_X1 _39579_ (.A(_14254_),
    .B(_14462_),
    .CI(_14463_),
    .CO(_14464_),
    .S(_14465_));
 FA_X1 _39580_ (.A(_14259_),
    .B(_14467_),
    .CI(_14466_),
    .CO(_14468_),
    .S(_14469_));
 FA_X1 _39581_ (.A(_14470_),
    .B(_14471_),
    .CI(_14468_),
    .CO(_14472_),
    .S(_14473_));
 FA_X1 _39582_ (.A(_14474_),
    .B(_14475_),
    .CI(_14476_),
    .CO(_14477_),
    .S(_14478_));
 FA_X1 _39583_ (.A(_14273_),
    .B(_14479_),
    .CI(_14480_),
    .CO(_14481_),
    .S(_14482_));
 FA_X1 _39584_ (.A(_14278_),
    .B(_14483_),
    .CI(_14484_),
    .CO(_14485_),
    .S(_14486_));
 FA_X1 _39585_ (.A(_14487_),
    .B(_14485_),
    .CI(_14488_),
    .CO(_14489_),
    .S(_14490_));
 FA_X1 _39586_ (.A(_14491_),
    .B(_14492_),
    .CI(_14493_),
    .CO(_14494_),
    .S(_14495_));
 FA_X1 _39587_ (.A(_14493_),
    .B(_14496_),
    .CI(_14497_),
    .CO(_14498_),
    .S(_14499_));
 FA_X1 _39588_ (.A(_14500_),
    .B(_14501_),
    .CI(_14502_),
    .CO(_14503_),
    .S(_14504_));
 FA_X1 _39589_ (.A(_14507_),
    .B(_14508_),
    .CI(_14509_),
    .CO(_14510_),
    .S(_14511_));
 FA_X1 _39590_ (.A(_14512_),
    .B(_14513_),
    .CI(_14509_),
    .CO(_14514_),
    .S(_14515_));
 FA_X1 _39591_ (.A(_14516_),
    .B(_14517_),
    .CI(_14518_),
    .CO(_14519_),
    .S(_14520_));
 FA_X1 _39592_ (.A(_14522_),
    .B(_14523_),
    .CI(_14524_),
    .CO(_14525_),
    .S(_14526_));
 FA_X1 _39593_ (.A(_14527_),
    .B(_14528_),
    .CI(_14529_),
    .CO(_14530_),
    .S(_14531_));
 FA_X1 _39594_ (.A(_14532_),
    .B(_14533_),
    .CI(_14534_),
    .CO(_14535_),
    .S(_14536_));
 FA_X1 _39595_ (.A(_14526_),
    .B(_14537_),
    .CI(_14538_),
    .CO(_14539_),
    .S(_14540_));
 FA_X1 _39596_ (.A(_14541_),
    .B(_14542_),
    .CI(_14543_),
    .CO(_14544_),
    .S(_14545_));
 FA_X1 _39597_ (.A(_14546_),
    .B(_14547_),
    .CI(_14548_),
    .CO(_14549_),
    .S(_14550_));
 FA_X1 _39598_ (.A(_14551_),
    .B(_14552_),
    .CI(_14553_),
    .CO(_14554_),
    .S(_14555_));
 FA_X1 _39599_ (.A(_14556_),
    .B(_14545_),
    .CI(_14557_),
    .CO(_14558_),
    .S(_14559_));
 FA_X1 _39600_ (.A(_14560_),
    .B(_14561_),
    .CI(_14562_),
    .CO(_14556_),
    .S(_14563_));
 FA_X1 _39601_ (.A(_14564_),
    .B(_14565_),
    .CI(_14566_),
    .CO(_14567_),
    .S(_14568_));
 FA_X1 _39602_ (.A(_14569_),
    .B(_14570_),
    .CI(_14571_),
    .CO(_14572_),
    .S(_14573_));
 FA_X1 _39603_ (.A(net266),
    .B(_14574_),
    .CI(_14575_),
    .CO(_14576_),
    .S(_14577_));
 FA_X1 _39604_ (.A(net83),
    .B(_14579_),
    .CI(_14580_),
    .CO(_14575_),
    .S(_14581_));
 FA_X1 _39605_ (.A(net82),
    .B(_14582_),
    .CI(_14583_),
    .CO(_14584_),
    .S(_14585_));
 FA_X1 _39606_ (.A(_14586_),
    .B(_14587_),
    .CI(_14588_),
    .CO(_14557_),
    .S(_14589_));
 FA_X1 _39607_ (.A(_14563_),
    .B(_14590_),
    .CI(_14591_),
    .CO(_14592_),
    .S(_14593_));
 FA_X1 _39608_ (.A(_14594_),
    .B(_14595_),
    .CI(_14596_),
    .CO(_14597_),
    .S(_14598_));
 FA_X1 _39609_ (.A(_14599_),
    .B(_14568_),
    .CI(_14600_),
    .CO(_14601_),
    .S(_14602_));
 FA_X1 _39610_ (.A(_14603_),
    .B(_14604_),
    .CI(_14605_),
    .CO(_14606_),
    .S(_14607_));
 FA_X1 _39611_ (.A(_14608_),
    .B(_14609_),
    .CI(_14610_),
    .CO(_14611_),
    .S(_14612_));
 FA_X1 _39612_ (.A(net84),
    .B(net267),
    .CI(_14613_),
    .CO(_14614_),
    .S(_14615_));
 FA_X1 _39613_ (.A(_14616_),
    .B(_14617_),
    .CI(_14618_),
    .CO(_14605_),
    .S(_14619_));
 FA_X1 _39614_ (.A(_14612_),
    .B(_14620_),
    .CI(_14621_),
    .CO(_14622_),
    .S(_14623_));
 FA_X1 _39615_ (.A(_14624_),
    .B(_14625_),
    .CI(_14626_),
    .CO(_14620_),
    .S(_14627_));
 FA_X1 _39616_ (.A(_14628_),
    .B(_14629_),
    .CI(_14630_),
    .CO(_14631_),
    .S(_14632_));
 FA_X1 _39617_ (.A(_14633_),
    .B(_14634_),
    .CI(_14635_),
    .CO(_14636_),
    .S(_14637_));
 FA_X1 _39618_ (.A(net61),
    .B(_14638_),
    .CI(_14639_),
    .CO(_14640_),
    .S(_14641_));
 FA_X1 _39619_ (.A(_14642_),
    .B(_14643_),
    .CI(_14644_),
    .CO(_14645_),
    .S(_14646_));
 FA_X1 _39620_ (.A(_14647_),
    .B(_14648_),
    .CI(_14649_),
    .CO(_14650_),
    .S(_14651_));
 FA_X1 _39621_ (.A(_14652_),
    .B(_14653_),
    .CI(_14654_),
    .CO(_14644_),
    .S(_14655_));
 FA_X1 _39622_ (.A(net250),
    .B(_14656_),
    .CI(_14657_),
    .CO(_14658_),
    .S(_14659_));
 FA_X1 _39623_ (.A(_14646_),
    .B(_14660_),
    .CI(_14661_),
    .CO(_14662_),
    .S(_14663_));
 FA_X1 _39624_ (.A(_14664_),
    .B(_14665_),
    .CI(_14666_),
    .CO(_14667_),
    .S(_14668_));
 FA_X1 _39625_ (.A(net62),
    .B(_14669_),
    .CI(_14670_),
    .CO(_14671_),
    .S(_14672_));
 FA_X1 _39626_ (.A(_14673_),
    .B(_14674_),
    .CI(_14672_),
    .CO(_14675_),
    .S(_14676_));
 FA_X1 _39627_ (.A(_14677_),
    .B(_14678_),
    .CI(_14679_),
    .CO(_14680_),
    .S(_14681_));
 FA_X1 _39628_ (.A(_14682_),
    .B(_14683_),
    .CI(_14681_),
    .CO(_14684_),
    .S(_14685_));
 FA_X1 _39629_ (.A(_14686_),
    .B(_14687_),
    .CI(_14688_),
    .CO(_14660_),
    .S(_14689_));
 FA_X1 _39630_ (.A(_14690_),
    .B(_14691_),
    .CI(_14692_),
    .CO(_14693_),
    .S(_14694_));
 FA_X1 _39631_ (.A(_14695_),
    .B(_14696_),
    .CI(_14697_),
    .CO(_14687_),
    .S(_14698_));
 FA_X1 _39632_ (.A(_14699_),
    .B(_14700_),
    .CI(_14701_),
    .CO(_14702_),
    .S(_14703_));
 FA_X1 _39633_ (.A(_14704_),
    .B(_14705_),
    .CI(_14706_),
    .CO(_14707_),
    .S(_14708_));
 FA_X1 _39634_ (.A(_14709_),
    .B(_14710_),
    .CI(_14711_),
    .CO(_14712_),
    .S(_14713_));
 FA_X1 _39635_ (.A(_14714_),
    .B(_14715_),
    .CI(_14716_),
    .CO(_14717_),
    .S(_14718_));
 FA_X1 _39636_ (.A(_14719_),
    .B(_14720_),
    .CI(_14721_),
    .CO(_14722_),
    .S(_14723_));
 FA_X1 _39637_ (.A(_14724_),
    .B(_14725_),
    .CI(_14726_),
    .CO(_14727_),
    .S(_14728_));
 FA_X1 _39638_ (.A(_14712_),
    .B(_14729_),
    .CI(_14728_),
    .CO(_14730_),
    .S(_14731_));
 FA_X1 _39639_ (.A(_14732_),
    .B(_14733_),
    .CI(_14734_),
    .CO(_14735_),
    .S(_14736_));
 FA_X1 _39640_ (.A(_14737_),
    .B(_14738_),
    .CI(_14736_),
    .CO(_14739_),
    .S(_14740_));
 FA_X1 _39641_ (.A(_14741_),
    .B(_14742_),
    .CI(_14743_),
    .CO(_14744_),
    .S(_14745_));
 FA_X1 _39642_ (.A(_14746_),
    .B(_14722_),
    .CI(_14747_),
    .CO(_14748_),
    .S(_14749_));
 FA_X1 _39643_ (.A(_14750_),
    .B(_14751_),
    .CI(_14752_),
    .CO(_14753_),
    .S(_14754_));
 FA_X1 _39644_ (.A(_14755_),
    .B(_14756_),
    .CI(_14757_),
    .CO(_14758_),
    .S(_14759_));
 FA_X1 _39645_ (.A(_14760_),
    .B(_14761_),
    .CI(_14762_),
    .CO(_14763_),
    .S(_14764_));
 FA_X1 _39646_ (.A(_14765_),
    .B(_14766_),
    .CI(_14767_),
    .CO(_14768_),
    .S(_14769_));
 FA_X1 _39647_ (.A(_14769_),
    .B(_14770_),
    .CI(_14771_),
    .CO(_14772_),
    .S(_14773_));
 FA_X1 _39648_ (.A(_14774_),
    .B(_14775_),
    .CI(_14776_),
    .CO(_14777_),
    .S(_14778_));
 FA_X1 _39649_ (.A(_14779_),
    .B(_14780_),
    .CI(_14781_),
    .CO(_14782_),
    .S(_14783_));
 FA_X1 _39650_ (.A(_14784_),
    .B(_14785_),
    .CI(_14786_),
    .CO(_14787_),
    .S(_14788_));
 FA_X1 _39651_ (.A(_14789_),
    .B(_14790_),
    .CI(_14783_),
    .CO(_14791_),
    .S(_14792_));
 FA_X1 _39652_ (.A(_14753_),
    .B(_14793_),
    .CI(_14758_),
    .CO(_14794_),
    .S(_14795_));
 FA_X1 _39653_ (.A(_14768_),
    .B(_14796_),
    .CI(_14763_),
    .CO(_14797_),
    .S(_14798_));
 FA_X1 _39654_ (.A(net141),
    .B(_14799_),
    .CI(_14800_),
    .CO(_14801_),
    .S(_14802_));
 FA_X1 _39655_ (.A(_14802_),
    .B(_14803_),
    .CI(_14804_),
    .CO(_14805_),
    .S(_14806_));
 FA_X1 _39656_ (.A(_14807_),
    .B(_14808_),
    .CI(_14809_),
    .CO(_14810_),
    .S(_14811_));
 FA_X1 _39657_ (.A(net261),
    .B(_14812_),
    .CI(_14813_),
    .CO(_14814_),
    .S(_14815_));
 FA_X1 _39658_ (.A(_14816_),
    .B(_14817_),
    .CI(_14818_),
    .CO(_14819_),
    .S(_14820_));
 FA_X1 _39659_ (.A(_14782_),
    .B(_14821_),
    .CI(_14822_),
    .CO(_14823_),
    .S(_14824_));
 FA_X1 _39660_ (.A(_14824_),
    .B(_14825_),
    .CI(_14791_),
    .CO(_14826_),
    .S(_14827_));
 FA_X1 _39661_ (.A(net142),
    .B(_14828_),
    .CI(_14829_),
    .CO(_14830_),
    .S(_14831_));
 FA_X1 _39662_ (.A(_14832_),
    .B(_14833_),
    .CI(_14831_),
    .CO(_14834_),
    .S(_14835_));
 FA_X1 _39663_ (.A(_14836_),
    .B(_14837_),
    .CI(_14838_),
    .CO(_14839_),
    .S(_14840_));
 FA_X1 _39664_ (.A(_14841_),
    .B(_14842_),
    .CI(_14843_),
    .CO(_14844_),
    .S(_14845_));
 FA_X1 _39665_ (.A(_14846_),
    .B(_14847_),
    .CI(_14845_),
    .CO(_14848_),
    .S(_14849_));
 FA_X1 _39666_ (.A(_14850_),
    .B(_14851_),
    .CI(_14852_),
    .CO(_14853_),
    .S(_14854_));
 FA_X1 _39667_ (.A(_14854_),
    .B(_14819_),
    .CI(_14823_),
    .CO(_14855_),
    .S(_14856_));
 FA_X1 _39668_ (.A(_14857_),
    .B(_14858_),
    .CI(_14859_),
    .CO(_14860_),
    .S(_14861_));
 FA_X1 _39669_ (.A(net143),
    .B(_14862_),
    .CI(_14863_),
    .CO(_14864_),
    .S(_14865_));
 FA_X1 _39670_ (.A(_14866_),
    .B(_14865_),
    .CI(_14830_),
    .CO(_14867_),
    .S(_14868_));
 FA_X1 _39671_ (.A(net263),
    .B(_14869_),
    .CI(_14870_),
    .CO(_14871_),
    .S(_14872_));
 FA_X1 _39672_ (.A(_14873_),
    .B(_14874_),
    .CI(_14875_),
    .CO(_14876_),
    .S(_14877_));
 FA_X1 _39673_ (.A(_14878_),
    .B(_14879_),
    .CI(_14844_),
    .CO(_14880_),
    .S(_14881_));
 FA_X1 _39674_ (.A(_14881_),
    .B(_14848_),
    .CI(_14853_),
    .CO(_14882_),
    .S(_14883_));
 FA_X1 _39675_ (.A(net144),
    .B(_14884_),
    .CI(_14885_),
    .CO(_14886_),
    .S(_14887_));
 FA_X1 _39676_ (.A(_14888_),
    .B(_14889_),
    .CI(_14890_),
    .CO(_14891_),
    .S(_14892_));
 FA_X1 _39677_ (.A(_14893_),
    .B(_14894_),
    .CI(_14895_),
    .CO(_14896_),
    .S(_14897_));
 FA_X1 _39678_ (.A(_14892_),
    .B(_14898_),
    .CI(_14899_),
    .CO(_14900_),
    .S(_14901_));
 FA_X1 _39679_ (.A(_14902_),
    .B(_14903_),
    .CI(_14904_),
    .CO(_14905_),
    .S(_14906_));
 FA_X1 _39680_ (.A(_14880_),
    .B(_14876_),
    .CI(_14906_),
    .CO(_14907_),
    .S(_14908_));
 FA_X1 _39681_ (.A(_14909_),
    .B(_14910_),
    .CI(_14911_),
    .CO(_14912_),
    .S(_14913_));
 FA_X1 _39682_ (.A(net145),
    .B(_14914_),
    .CI(_14915_),
    .CO(_14916_),
    .S(_14917_));
 FA_X1 _39683_ (.A(_14891_),
    .B(_14918_),
    .CI(_14919_),
    .CO(_14920_),
    .S(_14921_));
 FA_X1 _39684_ (.A(net264),
    .B(_14886_),
    .CI(_14896_),
    .CO(_14922_),
    .S(_14923_));
 FA_X1 _39685_ (.A(_14905_),
    .B(_14924_),
    .CI(_14900_),
    .CO(_14925_),
    .S(_14926_));
 FA_X1 _39686_ (.A(net146),
    .B(_14927_),
    .CI(_14928_),
    .CO(_14929_),
    .S(_14930_));
 FA_X1 _39687_ (.A(_14931_),
    .B(_14932_),
    .CI(_14933_),
    .CO(_14934_),
    .S(_14935_));
 FA_X1 _39688_ (.A(net265),
    .B(_14936_),
    .CI(_14937_),
    .CO(_14938_),
    .S(_14939_));
 FA_X1 _39689_ (.A(_14940_),
    .B(_14941_),
    .CI(_14920_),
    .CO(_14942_),
    .S(_14943_));
 FA_X1 _39690_ (.A(_14944_),
    .B(_14945_),
    .CI(_14946_),
    .CO(_14947_),
    .S(_14948_));
 FA_X1 _39691_ (.A(net147),
    .B(_14949_),
    .CI(_14950_),
    .CO(_14951_),
    .S(_14952_));
 FA_X1 _39692_ (.A(_14934_),
    .B(_14953_),
    .CI(_14954_),
    .CO(_14955_),
    .S(_14956_));
 FA_X1 _39693_ (.A(_14957_),
    .B(_14958_),
    .CI(_14959_),
    .CO(_14960_),
    .S(_14961_));
 FA_X1 _39694_ (.A(net266),
    .B(_14962_),
    .CI(_14951_),
    .CO(_14963_),
    .S(_14964_));
 FA_X1 _39695_ (.A(net148),
    .B(net267),
    .CI(_14965_),
    .CO(_14966_),
    .S(_14967_));
 FA_X1 _39696_ (.A(_14968_),
    .B(_14969_),
    .CI(_14970_),
    .CO(_14971_),
    .S(_14972_));
 FA_X1 _39697_ (.A(net28),
    .B(_14973_),
    .CI(_14974_),
    .CO(_14975_),
    .S(_14976_));
 FA_X1 _39698_ (.A(_14977_),
    .B(_14978_),
    .CI(_14976_),
    .CO(_14979_),
    .S(_14980_));
 FA_X1 _39699_ (.A(net232),
    .B(_14981_),
    .CI(_14982_),
    .CO(_14983_),
    .S(_14984_));
 FA_X1 _39700_ (.A(_14985_),
    .B(_14986_),
    .CI(_14987_),
    .CO(_14988_),
    .S(_14989_));
 FA_X1 _39701_ (.A(_14990_),
    .B(_14525_),
    .CI(_14991_),
    .CO(_14992_),
    .S(_14993_));
 FA_X1 _39702_ (.A(_14544_),
    .B(_14993_),
    .CI(_14539_),
    .CO(_14994_),
    .S(_14995_));
 FA_X1 _39703_ (.A(_14996_),
    .B(_14997_),
    .CI(_14998_),
    .CO(_14999_),
    .S(_15000_));
 FA_X1 _39704_ (.A(_15001_),
    .B(_15002_),
    .CI(_15003_),
    .CO(_14996_),
    .S(_15004_));
 FA_X1 _39705_ (.A(_15005_),
    .B(_15006_),
    .CI(_15007_),
    .CO(_14998_),
    .S(_15008_));
 FA_X1 _39706_ (.A(_15009_),
    .B(_15010_),
    .CI(_15011_),
    .CO(_15012_),
    .S(_15013_));
 FA_X1 _39707_ (.A(_15014_),
    .B(_15015_),
    .CI(_15016_),
    .CO(_15017_),
    .S(_15018_));
 FA_X1 _39708_ (.A(_15019_),
    .B(_15020_),
    .CI(_15021_),
    .CO(_15022_),
    .S(_15023_));
 FA_X1 _39709_ (.A(_15024_),
    .B(_15025_),
    .CI(_15026_),
    .CO(_15027_),
    .S(_15028_));
 FA_X1 _39710_ (.A(_15029_),
    .B(_15023_),
    .CI(_15030_),
    .CO(_15031_),
    .S(_15032_));
 FA_X1 _39711_ (.A(_15033_),
    .B(_15034_),
    .CI(_15035_),
    .CO(_15010_),
    .S(_15036_));
 FA_X1 _39712_ (.A(_15037_),
    .B(_15038_),
    .CI(_15039_),
    .CO(_15040_),
    .S(_15041_));
 FA_X1 _39713_ (.A(_15042_),
    .B(_15022_),
    .CI(_15043_),
    .CO(_15044_),
    .S(_15045_));
 FA_X1 _39714_ (.A(_15045_),
    .B(_15046_),
    .CI(_15031_),
    .CO(_15047_),
    .S(_15048_));
 FA_X1 _39715_ (.A(_15049_),
    .B(_15050_),
    .CI(_15051_),
    .CO(_15052_),
    .S(_15053_));
 FA_X1 _39716_ (.A(net76),
    .B(_15054_),
    .CI(_15055_),
    .CO(_15056_),
    .S(_15057_));
 FA_X1 _39717_ (.A(_15058_),
    .B(_15059_),
    .CI(_15060_),
    .CO(_15061_),
    .S(_15062_));
 FA_X1 _39718_ (.A(net261),
    .B(_15063_),
    .CI(_15064_),
    .CO(_15065_),
    .S(_15066_));
 FA_X1 _39719_ (.A(_15067_),
    .B(_15068_),
    .CI(_15062_),
    .CO(_15069_),
    .S(_15070_));
 FA_X1 _39720_ (.A(_15071_),
    .B(_15072_),
    .CI(_15061_),
    .CO(_15073_),
    .S(_15074_));
 FA_X1 _39721_ (.A(_15074_),
    .B(_15044_),
    .CI(_15069_),
    .CO(_15075_),
    .S(_15076_));
 FA_X1 _39722_ (.A(net77),
    .B(_15077_),
    .CI(_15078_),
    .CO(_15079_),
    .S(_15080_));
 FA_X1 _39723_ (.A(_15081_),
    .B(_15082_),
    .CI(_15080_),
    .CO(_15083_),
    .S(_15084_));
 FA_X1 _39724_ (.A(_15085_),
    .B(_15086_),
    .CI(_15087_),
    .CO(_15088_),
    .S(_15089_));
 FA_X1 _39725_ (.A(_14841_),
    .B(_15090_),
    .CI(_15091_),
    .CO(_15092_),
    .S(_15093_));
 FA_X1 _39726_ (.A(_15094_),
    .B(_15095_),
    .CI(_15093_),
    .CO(_15096_),
    .S(_15097_));
 FA_X1 _39727_ (.A(_15098_),
    .B(_15092_),
    .CI(_15099_),
    .CO(_15100_),
    .S(_15101_));
 FA_X1 _39728_ (.A(_15073_),
    .B(_15101_),
    .CI(_15096_),
    .CO(_15102_),
    .S(_15103_));
 FA_X1 _39729_ (.A(net78),
    .B(_15104_),
    .CI(_15105_),
    .CO(_15106_),
    .S(_15107_));
 FA_X1 _39730_ (.A(_15108_),
    .B(_15079_),
    .CI(_15107_),
    .CO(_15109_),
    .S(_15110_));
 FA_X1 _39731_ (.A(_15111_),
    .B(_15112_),
    .CI(_15113_),
    .CO(_15114_),
    .S(_15115_));
 FA_X1 _39732_ (.A(net263),
    .B(_15116_),
    .CI(_15117_),
    .CO(_15118_),
    .S(_15119_));
 FA_X1 _39733_ (.A(_15120_),
    .B(_15121_),
    .CI(_15122_),
    .CO(_15123_),
    .S(_15124_));
 FA_X1 _39734_ (.A(net36),
    .B(net275),
    .CI(_15125_),
    .CO(_15126_),
    .S(_15127_));
 FA_X1 _39735_ (.A(_15128_),
    .B(_14680_),
    .CI(_15129_),
    .CO(_15130_),
    .S(_15131_));
 FA_X1 _39736_ (.A(_15131_),
    .B(_14645_),
    .CI(_14684_),
    .CO(_15132_),
    .S(_15133_));
 FA_X1 _39737_ (.A(_15134_),
    .B(_15135_),
    .CI(_15136_),
    .CO(_15137_),
    .S(_15138_));
 FA_X1 _39738_ (.A(net63),
    .B(_15139_),
    .CI(_15140_),
    .CO(_15141_),
    .S(_15142_));
 FA_X1 _39739_ (.A(_15142_),
    .B(_14671_),
    .CI(_15143_),
    .CO(_15144_),
    .S(_15145_));
 FA_X1 _39740_ (.A(net251),
    .B(_15146_),
    .CI(_15147_),
    .CO(_15148_),
    .S(_15149_));
 FA_X1 _39741_ (.A(_15150_),
    .B(_15151_),
    .CI(_15152_),
    .CO(_15153_),
    .S(_15154_));
 FA_X1 _39742_ (.A(_15155_),
    .B(_15156_),
    .CI(_15157_),
    .CO(_15158_),
    .S(_15159_));
 FA_X1 _39743_ (.A(net274),
    .B(_15160_),
    .CI(_15161_),
    .CO(_15162_),
    .S(_15163_));
 FA_X1 _39744_ (.A(net35),
    .B(_15165_),
    .CI(_15166_),
    .CO(_15160_),
    .S(_15167_));
 FA_X1 _39745_ (.A(net34),
    .B(_15168_),
    .CI(_15169_),
    .CO(_15170_),
    .S(_15171_));
 FA_X1 _39746_ (.A(net79),
    .B(_15172_),
    .CI(_15173_),
    .CO(_15174_),
    .S(_15175_));
 FA_X1 _39747_ (.A(_14888_),
    .B(_15176_),
    .CI(_15177_),
    .CO(_15178_),
    .S(_15179_));
 FA_X1 _39748_ (.A(_15180_),
    .B(_15181_),
    .CI(_15182_),
    .CO(_15183_),
    .S(_15184_));
 FA_X1 _39749_ (.A(_15185_),
    .B(_15179_),
    .CI(_15186_),
    .CO(_15187_),
    .S(_15188_));
 FA_X1 _39750_ (.A(_15189_),
    .B(_15190_),
    .CI(_15191_),
    .CO(_15192_),
    .S(_15193_));
 FA_X1 _39751_ (.A(_15100_),
    .B(_15193_),
    .CI(_15123_),
    .CO(_15194_),
    .S(_15195_));
 FA_X1 _39752_ (.A(_15196_),
    .B(_15197_),
    .CI(_15198_),
    .CO(_15164_),
    .S(_15199_));
 FA_X1 _39753_ (.A(_15200_),
    .B(_15201_),
    .CI(_15202_),
    .CO(_15203_),
    .S(_15204_));
 FA_X1 _39754_ (.A(net270),
    .B(_15205_),
    .CI(_15206_),
    .CO(_15207_),
    .S(_15208_));
 FA_X1 _39755_ (.A(_15209_),
    .B(_15210_),
    .CI(_15211_),
    .CO(_15212_),
    .S(_15213_));
 FA_X1 _39756_ (.A(net33),
    .B(_15214_),
    .CI(_15215_),
    .CO(_15216_),
    .S(_15217_));
 FA_X1 _39757_ (.A(_15218_),
    .B(_15219_),
    .CI(_15220_),
    .CO(_15202_),
    .S(_15221_));
 FA_X1 _39758_ (.A(_15222_),
    .B(_15223_),
    .CI(_15224_),
    .CO(_15225_),
    .S(_15226_));
 FA_X1 _39759_ (.A(net31),
    .B(_15227_),
    .CI(_15228_),
    .CO(_15229_),
    .S(_15230_));
 FA_X1 _39760_ (.A(net262),
    .B(_15231_),
    .CI(_15232_),
    .CO(_15233_),
    .S(_15234_));
 FA_X1 _39761_ (.A(net32),
    .B(_15235_),
    .CI(_15236_),
    .CO(_15232_),
    .S(_15237_));
 FA_X1 _39762_ (.A(_15238_),
    .B(_15239_),
    .CI(_15240_),
    .CO(_15241_),
    .S(_15242_));
 FA_X1 _39763_ (.A(_15243_),
    .B(_15244_),
    .CI(_15245_),
    .CO(_15231_),
    .S(_15246_));
 FA_X1 _39764_ (.A(_15247_),
    .B(_15248_),
    .CI(_15249_),
    .CO(_15250_),
    .S(_15251_));
 FA_X1 _39765_ (.A(net81),
    .B(_15252_),
    .CI(_15253_),
    .CO(_15254_),
    .S(_15255_));
 FA_X1 _39766_ (.A(_15256_),
    .B(_15178_),
    .CI(_15257_),
    .CO(_15258_),
    .S(_15259_));
 FA_X1 _39767_ (.A(net264),
    .B(_15174_),
    .CI(_15183_),
    .CO(_15260_),
    .S(_15261_));
 FA_X1 _39768_ (.A(_15262_),
    .B(_15192_),
    .CI(_15187_),
    .CO(_15263_),
    .S(_15264_));
 FA_X1 _39769_ (.A(_15265_),
    .B(_15241_),
    .CI(_15266_),
    .CO(_15224_),
    .S(_15267_));
 FA_X1 _39770_ (.A(_15268_),
    .B(_15269_),
    .CI(_15270_),
    .CO(_15271_),
    .S(_15272_));
 FA_X1 _39771_ (.A(_15273_),
    .B(_15274_),
    .CI(_15275_),
    .CO(_15268_),
    .S(_15276_));
 FA_X1 _39772_ (.A(net29),
    .B(_15277_),
    .CI(_15278_),
    .CO(_15279_),
    .S(_15280_));
 FA_X1 _39773_ (.A(_15281_),
    .B(_15282_),
    .CI(_15283_),
    .CO(_15284_),
    .S(_15285_));
 FA_X1 _39774_ (.A(_15279_),
    .B(_15230_),
    .CI(_15286_),
    .CO(_15287_),
    .S(_15288_));
 FA_X1 _39775_ (.A(net248),
    .B(_15289_),
    .CI(_15290_),
    .CO(_15291_),
    .S(_15292_));
 FA_X1 _39776_ (.A(_15293_),
    .B(_15242_),
    .CI(_15294_),
    .CO(_15270_),
    .S(_15295_));
 FA_X1 _39777_ (.A(_15276_),
    .B(_15296_),
    .CI(_15297_),
    .CO(_15298_),
    .S(_15299_));
 FA_X1 _39778_ (.A(_15300_),
    .B(_15301_),
    .CI(_15302_),
    .CO(_15296_),
    .S(_15303_));
 FA_X1 _39779_ (.A(_15304_),
    .B(_15305_),
    .CI(_15306_),
    .CO(_15307_),
    .S(_15308_));
 FA_X1 _39780_ (.A(_15309_),
    .B(_15310_),
    .CI(_15311_),
    .CO(_15300_),
    .S(_15312_));
 FA_X1 _39781_ (.A(_15313_),
    .B(_15314_),
    .CI(_15315_),
    .CO(_15302_),
    .S(_15316_));
 FA_X1 _39782_ (.A(_15317_),
    .B(_15318_),
    .CI(_15319_),
    .CO(_15320_),
    .S(_15321_));
 FA_X1 _39783_ (.A(net265),
    .B(_15322_),
    .CI(_15323_),
    .CO(_15324_),
    .S(_15325_));
 FA_X1 _39784_ (.A(_15326_),
    .B(_15327_),
    .CI(_15258_),
    .CO(_15328_),
    .S(_15329_));
 FA_X1 _39785_ (.A(_15330_),
    .B(_15331_),
    .CI(_15332_),
    .CO(_15297_),
    .S(_15333_));
 FA_X1 _39786_ (.A(_15303_),
    .B(_15334_),
    .CI(_15335_),
    .CO(_15336_),
    .S(_15337_));
 FA_X1 _39787_ (.A(_15338_),
    .B(_15339_),
    .CI(_15340_),
    .CO(_15334_),
    .S(_15341_));
 FA_X1 _39788_ (.A(_15312_),
    .B(_15342_),
    .CI(_15316_),
    .CO(_15335_),
    .S(_15343_));
 FA_X1 _39789_ (.A(_15341_),
    .B(_14992_),
    .CI(_14988_),
    .CO(_15344_),
    .S(_15345_));
 FA_X1 _39790_ (.A(_14944_),
    .B(_15346_),
    .CI(_15347_),
    .CO(_14578_),
    .S(_15348_));
 FA_X1 _39791_ (.A(_15349_),
    .B(_15350_),
    .CI(_15320_),
    .CO(_15351_),
    .S(_15352_));
 FA_X1 _39792_ (.A(_15353_),
    .B(_15354_),
    .CI(_15355_),
    .CO(_15356_),
    .S(_15357_));
 FA_X1 _39793_ (.A(_15358_),
    .B(_15359_),
    .CI(_15360_),
    .CO(_15361_),
    .S(_15362_));
 FA_X1 _39794_ (.A(_15363_),
    .B(_15364_),
    .CI(_15365_),
    .CO(_15366_),
    .S(_15367_));
 FA_X1 _39795_ (.A(_15368_),
    .B(_15369_),
    .CI(_15370_),
    .CO(_15371_),
    .S(_15372_));
 FA_X1 _39796_ (.A(_15373_),
    .B(_15374_),
    .CI(_15375_),
    .CO(_15376_),
    .S(_15377_));
 FA_X1 _39797_ (.A(_15377_),
    .B(_15361_),
    .CI(_15378_),
    .CO(_15379_),
    .S(_15380_));
 FA_X1 _39798_ (.A(_15381_),
    .B(_15382_),
    .CI(_15383_),
    .CO(_15384_),
    .S(_15385_));
 FA_X1 _39799_ (.A(_15386_),
    .B(_15387_),
    .CI(_15388_),
    .CO(_15389_),
    .S(_15390_));
 FA_X1 _39800_ (.A(_15384_),
    .B(_15391_),
    .CI(_15392_),
    .CO(_15393_),
    .S(_15394_));
 FA_X1 _39801_ (.A(_15395_),
    .B(_15396_),
    .CI(_15397_),
    .CO(_15398_),
    .S(_15399_));
 FA_X1 _39802_ (.A(_15400_),
    .B(_15401_),
    .CI(_15402_),
    .CO(_15403_),
    .S(_15404_));
 FA_X1 _39803_ (.A(_15405_),
    .B(_15406_),
    .CI(_15407_),
    .CO(_15408_),
    .S(_15409_));
 FA_X1 _39804_ (.A(_15130_),
    .B(_15409_),
    .CI(_15153_),
    .CO(_15410_),
    .S(_15411_));
 FA_X1 _39805_ (.A(_15412_),
    .B(_15413_),
    .CI(_15414_),
    .CO(_15415_),
    .S(_15416_));
 FA_X1 _39806_ (.A(net64),
    .B(_15417_),
    .CI(_15418_),
    .CO(_15419_),
    .S(_15420_));
 FA_X1 _39807_ (.A(_15421_),
    .B(_15422_),
    .CI(_15423_),
    .CO(_15424_),
    .S(_15425_));
 FA_X1 _39808_ (.A(_15426_),
    .B(_15416_),
    .CI(_15427_),
    .CO(_15428_),
    .S(_15429_));
 FA_X1 _39809_ (.A(_15430_),
    .B(_15431_),
    .CI(_15432_),
    .CO(_15433_),
    .S(_15434_));
 FA_X1 _39810_ (.A(_15435_),
    .B(_15434_),
    .CI(_15403_),
    .CO(_15436_),
    .S(_15437_));
 FA_X1 _39811_ (.A(_15438_),
    .B(_15439_),
    .CI(_15440_),
    .CO(_15441_),
    .S(_15442_));
 FA_X1 _39812_ (.A(_15443_),
    .B(_15444_),
    .CI(_15445_),
    .CO(_15446_),
    .S(_15447_));
 FA_X1 _39813_ (.A(_15448_),
    .B(_15449_),
    .CI(_15450_),
    .CO(_15451_),
    .S(_15452_));
 FA_X1 _39814_ (.A(_15453_),
    .B(_15441_),
    .CI(_15446_),
    .CO(_15454_),
    .S(_15455_));
 FA_X1 _39815_ (.A(_15456_),
    .B(_15433_),
    .CI(_15451_),
    .CO(_15457_),
    .S(_15458_));
 FA_X1 _39816_ (.A(_15459_),
    .B(_15460_),
    .CI(_15461_),
    .CO(_15462_),
    .S(_15463_));
 FA_X1 _39817_ (.A(_15464_),
    .B(_15465_),
    .CI(_15466_),
    .CO(_15467_),
    .S(_15468_));
 FA_X1 _39818_ (.A(_15469_),
    .B(_15470_),
    .CI(_15471_),
    .CO(_15472_),
    .S(_15473_));
 FA_X1 _39819_ (.A(_15474_),
    .B(_15463_),
    .CI(_15475_),
    .CO(_15476_),
    .S(_15477_));
 FA_X1 _39820_ (.A(_15478_),
    .B(_15479_),
    .CI(_15480_),
    .CO(_15481_),
    .S(_15482_));
 FA_X1 _39821_ (.A(_15483_),
    .B(_15484_),
    .CI(_15485_),
    .CO(_15486_),
    .S(_15487_));
 FA_X1 _39822_ (.A(_15462_),
    .B(_15488_),
    .CI(_15489_),
    .CO(_15490_),
    .S(_15491_));
 FA_X1 _39823_ (.A(_15491_),
    .B(_15492_),
    .CI(_15476_),
    .CO(_15493_),
    .S(_15494_));
 FA_X1 _39824_ (.A(_15495_),
    .B(_15496_),
    .CI(_15497_),
    .CO(_15498_),
    .S(_15499_));
 FA_X1 _39825_ (.A(net125),
    .B(_15500_),
    .CI(_15501_),
    .CO(_15502_),
    .S(_15503_));
 FA_X1 _39826_ (.A(_15504_),
    .B(_15505_),
    .CI(_15506_),
    .CO(_15507_),
    .S(_15508_));
 FA_X1 _39827_ (.A(net250),
    .B(_15509_),
    .CI(_15510_),
    .CO(_15511_),
    .S(_15512_));
 FA_X1 _39828_ (.A(_15513_),
    .B(_15508_),
    .CI(_15514_),
    .CO(_15515_),
    .S(_15516_));
 FA_X1 _39829_ (.A(_15517_),
    .B(_15507_),
    .CI(_15518_),
    .CO(_15519_),
    .S(_15520_));
 FA_X1 _39830_ (.A(_15520_),
    .B(_15490_),
    .CI(_15515_),
    .CO(_15521_),
    .S(_15522_));
 FA_X1 _39831_ (.A(_15523_),
    .B(_15524_),
    .CI(_15525_),
    .CO(_15526_),
    .S(_15527_));
 FA_X1 _39832_ (.A(net126),
    .B(_15528_),
    .CI(_15529_),
    .CO(_15530_),
    .S(_15531_));
 FA_X1 _39833_ (.A(_15532_),
    .B(_15533_),
    .CI(_15531_),
    .CO(_15534_),
    .S(_15535_));
 FA_X1 _39834_ (.A(_14677_),
    .B(_15536_),
    .CI(_15537_),
    .CO(_15538_),
    .S(_15539_));
 FA_X1 _39835_ (.A(_15540_),
    .B(_15541_),
    .CI(_15539_),
    .CO(_15542_),
    .S(_15543_));
 FA_X1 _39836_ (.A(_15544_),
    .B(_15545_),
    .CI(_15538_),
    .CO(_15546_),
    .S(_15547_));
 FA_X1 _39837_ (.A(_15547_),
    .B(_15542_),
    .CI(_15519_),
    .CO(_15548_),
    .S(_15549_));
 FA_X1 _39838_ (.A(_15550_),
    .B(_15551_),
    .CI(_15552_),
    .CO(_15553_),
    .S(_15554_));
 FA_X1 _39839_ (.A(net127),
    .B(_15555_),
    .CI(_15556_),
    .CO(_15557_),
    .S(_15558_));
 FA_X1 _39840_ (.A(_15558_),
    .B(_15559_),
    .CI(_15530_),
    .CO(_15560_),
    .S(_15561_));
 FA_X1 _39841_ (.A(net251),
    .B(_15562_),
    .CI(_15563_),
    .CO(_15564_),
    .S(_15565_));
 FA_X1 _39842_ (.A(_15566_),
    .B(_15567_),
    .CI(_15568_),
    .CO(_15569_),
    .S(_15570_));
 FA_X1 _39843_ (.A(_15571_),
    .B(_15572_),
    .CI(_15573_),
    .CO(_15574_),
    .S(_15575_));
 FA_X1 _39844_ (.A(_15575_),
    .B(_15546_),
    .CI(_15569_),
    .CO(_15576_),
    .S(_15577_));
 FA_X1 _39845_ (.A(_15412_),
    .B(_15578_),
    .CI(_15579_),
    .CO(_15580_),
    .S(_15581_));
 FA_X1 _39846_ (.A(net128),
    .B(_15582_),
    .CI(_15583_),
    .CO(_15584_),
    .S(_15585_));
 FA_X1 _39847_ (.A(_15586_),
    .B(_15587_),
    .CI(_15588_),
    .CO(_15589_),
    .S(_15590_));
 FA_X1 _39848_ (.A(_15581_),
    .B(_15591_),
    .CI(_15592_),
    .CO(_15593_),
    .S(_15594_));
 FA_X1 _39849_ (.A(_15595_),
    .B(_15596_),
    .CI(_15597_),
    .CO(_15598_),
    .S(_15599_));
 FA_X1 _39850_ (.A(_15481_),
    .B(_15600_),
    .CI(_15599_),
    .CO(_15601_),
    .S(_15602_));
 FA_X1 _39851_ (.A(_15603_),
    .B(_15604_),
    .CI(_15605_),
    .CO(_15606_),
    .S(_15607_));
 FA_X1 _39852_ (.A(net252),
    .B(_15584_),
    .CI(_15589_),
    .CO(_15608_),
    .S(_15609_));
 FA_X1 _39853_ (.A(_15610_),
    .B(_15574_),
    .CI(_15593_),
    .CO(_15611_),
    .S(_15612_));
 FA_X1 _39854_ (.A(_15613_),
    .B(_15614_),
    .CI(_15615_),
    .CO(_15616_),
    .S(_15617_));
 FA_X1 _39855_ (.A(net129),
    .B(_15618_),
    .CI(_15619_),
    .CO(_15620_),
    .S(_15621_));
 FA_X1 _39856_ (.A(_15580_),
    .B(_15622_),
    .CI(_15623_),
    .CO(_15624_),
    .S(_15625_));
 FA_X1 _39857_ (.A(net253),
    .B(_15626_),
    .CI(_15627_),
    .CO(_15628_),
    .S(_15629_));
 FA_X1 _39858_ (.A(_15630_),
    .B(_15624_),
    .CI(_15631_),
    .CO(_15632_),
    .S(_15633_));
 FA_X1 _39859_ (.A(net130),
    .B(_15634_),
    .CI(_15635_),
    .CO(_15636_),
    .S(_15637_));
 FA_X1 _39860_ (.A(_15638_),
    .B(_15639_),
    .CI(_15640_),
    .CO(_15641_),
    .S(_15642_));
 FA_X1 _39861_ (.A(net132),
    .B(_15643_),
    .CI(_15644_),
    .CO(_15645_),
    .S(_15646_));
 FA_X1 _39862_ (.A(_15647_),
    .B(_15648_),
    .CI(_15641_),
    .CO(_15649_),
    .S(_15650_));
 FA_X1 _39863_ (.A(_15651_),
    .B(_15652_),
    .CI(_15653_),
    .CO(_15654_),
    .S(_15655_));
 FA_X1 _39864_ (.A(net254),
    .B(_15645_),
    .CI(_15656_),
    .CO(_15657_),
    .S(_15658_));
 FA_X1 _39865_ (.A(net133),
    .B(_15659_),
    .CI(_15660_),
    .CO(_15661_),
    .S(_15662_));
 FA_X1 _39866_ (.A(_15663_),
    .B(_15664_),
    .CI(_15665_),
    .CO(_15666_),
    .S(_15667_));
 FA_X1 _39867_ (.A(_15668_),
    .B(_15669_),
    .CI(_15606_),
    .CO(_15670_),
    .S(_15671_));
 FA_X1 _39868_ (.A(_15672_),
    .B(_15673_),
    .CI(_15674_),
    .CO(_15675_),
    .S(_15676_));
 FA_X1 _39869_ (.A(net134),
    .B(net255),
    .CI(_15677_),
    .CO(_15678_),
    .S(_15679_));
 FA_X1 _39870_ (.A(_15675_),
    .B(_15680_),
    .CI(_15036_),
    .CO(_15681_),
    .S(_15682_));
 FA_X1 _39871_ (.A(_15683_),
    .B(_15684_),
    .CI(_15685_),
    .CO(_15011_),
    .S(_15686_));
 FA_X1 _39872_ (.A(_15687_),
    .B(_15688_),
    .CI(_15689_),
    .CO(_15690_),
    .S(_15691_));
 FA_X1 _39873_ (.A(net65),
    .B(_15692_),
    .CI(_15693_),
    .CO(_15694_),
    .S(_15695_));
 FA_X1 _39874_ (.A(_15696_),
    .B(_15415_),
    .CI(_15697_),
    .CO(_15698_),
    .S(_15699_));
 FA_X1 _39875_ (.A(net252),
    .B(_15424_),
    .CI(_15419_),
    .CO(_15700_),
    .S(_15701_));
 FA_X1 _39876_ (.A(_15408_),
    .B(_15702_),
    .CI(_15428_),
    .CO(_15703_),
    .S(_15704_));
 FA_X1 _39877_ (.A(net68),
    .B(net255),
    .CI(_15705_),
    .CO(_15706_),
    .S(_15707_));
 FA_X1 _39878_ (.A(_15708_),
    .B(_15709_),
    .CI(_15710_),
    .CO(_15711_),
    .S(_15712_));
 FA_X1 _39879_ (.A(_15713_),
    .B(_15714_),
    .CI(_15715_),
    .CO(_15716_),
    .S(_15717_));
 FA_X1 _39880_ (.A(_15718_),
    .B(_15719_),
    .CI(_15720_),
    .CO(_15721_),
    .S(_15722_));
 FA_X1 _39881_ (.A(_15723_),
    .B(_15724_),
    .CI(_15725_),
    .CO(_15726_),
    .S(_15727_));
 FA_X1 _39882_ (.A(_15716_),
    .B(_15728_),
    .CI(_15727_),
    .CO(_15729_),
    .S(_15730_));
 FA_X1 _39883_ (.A(_15731_),
    .B(_15732_),
    .CI(_15733_),
    .CO(_15734_),
    .S(_15735_));
 FA_X1 _39884_ (.A(_15736_),
    .B(_15737_),
    .CI(_15738_),
    .CO(_15739_),
    .S(_15740_));
 FA_X1 _39885_ (.A(_15741_),
    .B(_15742_),
    .CI(_15734_),
    .CO(_15743_),
    .S(_15744_));
 FA_X1 _39886_ (.A(_15745_),
    .B(_15746_),
    .CI(_15747_),
    .CO(_15748_),
    .S(_15749_));
 FA_X1 _39887_ (.A(_15750_),
    .B(_15751_),
    .CI(_15749_),
    .CO(_15752_),
    .S(_15753_));
 FA_X1 _39888_ (.A(net66),
    .B(_15754_),
    .CI(_15755_),
    .CO(_15756_),
    .S(_15757_));
 FA_X1 _39889_ (.A(_15758_),
    .B(_15759_),
    .CI(_15760_),
    .CO(_15761_),
    .S(_15762_));
 FA_X1 _39890_ (.A(net253),
    .B(_15763_),
    .CI(_15764_),
    .CO(_15765_),
    .S(_15766_));
 FA_X1 _39891_ (.A(_15698_),
    .B(_15767_),
    .CI(_15768_),
    .CO(_15769_),
    .S(_15770_));
 FA_X1 _39892_ (.A(_15771_),
    .B(_15772_),
    .CI(_15773_),
    .CO(_15774_),
    .S(_15775_));
 FA_X1 _39893_ (.A(_15776_),
    .B(_15777_),
    .CI(_15775_),
    .CO(_15778_),
    .S(_15779_));
 FA_X1 _39894_ (.A(_15780_),
    .B(_15781_),
    .CI(_15782_),
    .CO(_15783_),
    .S(_15784_));
 FA_X1 _39895_ (.A(_15785_),
    .B(_15786_),
    .CI(_15787_),
    .CO(_15788_),
    .S(_15789_));
 FA_X1 _39896_ (.A(_15790_),
    .B(_15791_),
    .CI(_15792_),
    .CO(_15793_),
    .S(_15794_));
 FA_X1 _39897_ (.A(_15788_),
    .B(_15783_),
    .CI(_15795_),
    .CO(_15796_),
    .S(_15797_));
 FA_X1 _39898_ (.A(_15798_),
    .B(_15774_),
    .CI(_15793_),
    .CO(_15799_),
    .S(_15800_));
 FA_X1 _39899_ (.A(_15801_),
    .B(_15802_),
    .CI(_15803_),
    .CO(_15804_),
    .S(_15805_));
 FA_X1 _39900_ (.A(_15806_),
    .B(_15807_),
    .CI(_15808_),
    .CO(_15809_),
    .S(_15810_));
 FA_X1 _39901_ (.A(_15811_),
    .B(_15812_),
    .CI(_15813_),
    .CO(_15814_),
    .S(_15815_));
 FA_X1 _39902_ (.A(_15816_),
    .B(_15810_),
    .CI(_15817_),
    .CO(_15818_),
    .S(_15819_));
 FA_X1 _39903_ (.A(_15809_),
    .B(_15820_),
    .CI(_15821_),
    .CO(_15822_),
    .S(_15823_));
 FA_X1 _39904_ (.A(_15823_),
    .B(_15824_),
    .CI(_15818_),
    .CO(_15825_),
    .S(_15826_));
 FA_X1 _39905_ (.A(net108),
    .B(_15827_),
    .CI(_15828_),
    .CO(_15829_),
    .S(_15830_));
 FA_X1 _39906_ (.A(_15831_),
    .B(_15832_),
    .CI(_15830_),
    .CO(_15833_),
    .S(_15834_));
 FA_X1 _39907_ (.A(_15835_),
    .B(_15836_),
    .CI(_15837_),
    .CO(_15838_),
    .S(_15839_));
 FA_X1 _39908_ (.A(net238),
    .B(_15840_),
    .CI(_15841_),
    .CO(_15842_),
    .S(_15843_));
 FA_X1 _39909_ (.A(_15844_),
    .B(_15845_),
    .CI(_15846_),
    .CO(_15847_),
    .S(_15848_));
 FA_X1 _39910_ (.A(_15849_),
    .B(_15850_),
    .CI(_15851_),
    .CO(_15852_),
    .S(_15853_));
 FA_X1 _39911_ (.A(_15853_),
    .B(_15822_),
    .CI(_15847_),
    .CO(_15854_),
    .S(_15855_));
 FA_X1 _39912_ (.A(_15856_),
    .B(_15857_),
    .CI(_15858_),
    .CO(_15859_),
    .S(_15860_));
 FA_X1 _39913_ (.A(net109),
    .B(_15861_),
    .CI(_15862_),
    .CO(_15863_),
    .S(_15864_));
 FA_X1 _39914_ (.A(_15865_),
    .B(_15866_),
    .CI(_15867_),
    .CO(_15868_),
    .S(_15869_));
 FA_X1 _39915_ (.A(_15870_),
    .B(_15871_),
    .CI(_15872_),
    .CO(_15873_),
    .S(_15874_));
 FA_X1 _39916_ (.A(_15874_),
    .B(_15875_),
    .CI(_15869_),
    .CO(_15876_),
    .S(_15877_));
 FA_X1 _39917_ (.A(_15868_),
    .B(_15878_),
    .CI(_15873_),
    .CO(_15879_),
    .S(_15880_));
 FA_X1 _39918_ (.A(_15880_),
    .B(_15852_),
    .CI(_15876_),
    .CO(_15881_),
    .S(_15882_));
 FA_X1 _39919_ (.A(net111),
    .B(_15883_),
    .CI(_15884_),
    .CO(_15885_),
    .S(_15886_));
 FA_X1 _39920_ (.A(_15886_),
    .B(_15863_),
    .CI(_15887_),
    .CO(_15888_),
    .S(_15889_));
 FA_X1 _39921_ (.A(_15890_),
    .B(_15891_),
    .CI(_15892_),
    .CO(_15893_),
    .S(_15894_));
 FA_X1 _39922_ (.A(net239),
    .B(_15895_),
    .CI(_15896_),
    .CO(_15897_),
    .S(_15898_));
 FA_X1 _39923_ (.A(_15899_),
    .B(_15900_),
    .CI(_15901_),
    .CO(_15902_),
    .S(_15903_));
 FA_X1 _39924_ (.A(_15904_),
    .B(_15905_),
    .CI(_15906_),
    .CO(_15907_),
    .S(_15908_));
 FA_X1 _39925_ (.A(_15879_),
    .B(_15902_),
    .CI(_15908_),
    .CO(_15909_),
    .S(_15910_));
 FA_X1 _39926_ (.A(net112),
    .B(_15911_),
    .CI(_15912_),
    .CO(_15913_),
    .S(_15914_));
 FA_X1 _39927_ (.A(_15915_),
    .B(_15916_),
    .CI(_15917_),
    .CO(_15918_),
    .S(_15919_));
 FA_X1 _39928_ (.A(_15920_),
    .B(_15921_),
    .CI(_15922_),
    .CO(_15923_),
    .S(_15924_));
 FA_X1 _39929_ (.A(_15925_),
    .B(_15919_),
    .CI(_15926_),
    .CO(_15927_),
    .S(_15928_));
 FA_X1 _39930_ (.A(_15929_),
    .B(_15930_),
    .CI(_15931_),
    .CO(_15932_),
    .S(_15933_));
 FA_X1 _39931_ (.A(net113),
    .B(_15934_),
    .CI(_15935_),
    .CO(_15936_),
    .S(_15937_));
 FA_X1 _39932_ (.A(_15938_),
    .B(_15918_),
    .CI(_15939_),
    .CO(_15940_),
    .S(_15941_));
 FA_X1 _39933_ (.A(net240),
    .B(_15923_),
    .CI(_15913_),
    .CO(_15942_),
    .S(_15943_));
 FA_X1 _39934_ (.A(_15944_),
    .B(_15907_),
    .CI(_15927_),
    .CO(_15945_),
    .S(_15946_));
 FA_X1 _39935_ (.A(net114),
    .B(_15947_),
    .CI(_15948_),
    .CO(_15949_),
    .S(_15950_));
 FA_X1 _39936_ (.A(_15951_),
    .B(_15952_),
    .CI(_15953_),
    .CO(_15954_),
    .S(_15955_));
 FA_X1 _39937_ (.A(net241),
    .B(_15956_),
    .CI(_15957_),
    .CO(_15958_),
    .S(_15959_));
 FA_X1 _39938_ (.A(_15940_),
    .B(_15960_),
    .CI(_15961_),
    .CO(_15962_),
    .S(_15963_));
 FA_X1 _39939_ (.A(_15964_),
    .B(_15965_),
    .CI(_15966_),
    .CO(_15967_),
    .S(_15968_));
 FA_X1 _39940_ (.A(net115),
    .B(_15969_),
    .CI(_15970_),
    .CO(_15971_),
    .S(_15972_));
 FA_X1 _39941_ (.A(_15973_),
    .B(_15974_),
    .CI(_15954_),
    .CO(_15975_),
    .S(_15976_));
 FA_X1 _39942_ (.A(net242),
    .B(_15977_),
    .CI(_15971_),
    .CO(_15978_),
    .S(_15979_));
 FA_X1 _39943_ (.A(net116),
    .B(_15980_),
    .CI(_15981_),
    .CO(_15982_),
    .S(_15983_));
 FA_X1 _39944_ (.A(net117),
    .B(net243),
    .CI(_15984_),
    .CO(_15985_),
    .S(_15986_));
 FA_X1 _39945_ (.A(net241),
    .B(_15987_),
    .CI(_15988_),
    .CO(_15989_),
    .S(_15990_));
 FA_X1 _39946_ (.A(_15991_),
    .B(_15992_),
    .CI(_15993_),
    .CO(_15994_),
    .S(_15995_));
 FA_X1 _39947_ (.A(net48),
    .B(_15996_),
    .CI(_15997_),
    .CO(_15998_),
    .S(_15999_));
 FA_X1 _39948_ (.A(_16000_),
    .B(_16001_),
    .CI(_16002_),
    .CO(_16003_),
    .S(_16004_));
 FA_X1 _39949_ (.A(net49),
    .B(_16005_),
    .CI(_16006_),
    .CO(_16007_),
    .S(_16008_));
 FA_X1 _39950_ (.A(_16009_),
    .B(_16010_),
    .CI(_16011_),
    .CO(_16012_),
    .S(_16013_));
 FA_X1 _39951_ (.A(net240),
    .B(_16014_),
    .CI(_16015_),
    .CO(_16016_),
    .S(_16017_));
 FA_X1 _39952_ (.A(net46),
    .B(_16018_),
    .CI(_16019_),
    .CO(_16020_),
    .S(_16021_));
 FA_X1 _39953_ (.A(net47),
    .B(_16022_),
    .CI(_16023_),
    .CO(_16015_),
    .S(_16024_));
 FA_X1 _39954_ (.A(_15915_),
    .B(_16025_),
    .CI(_16026_),
    .CO(_16027_),
    .S(_16028_));
 FA_X1 _39955_ (.A(_16029_),
    .B(_16030_),
    .CI(_16031_),
    .CO(_16014_),
    .S(_16032_));
 FA_X1 _39956_ (.A(_16033_),
    .B(_16034_),
    .CI(_16035_),
    .CO(_16036_),
    .S(_16037_));
 FA_X1 _39957_ (.A(_16038_),
    .B(_16027_),
    .CI(_16039_),
    .CO(_16002_),
    .S(_16040_));
 FA_X1 _39958_ (.A(net45),
    .B(_16041_),
    .CI(_16042_),
    .CO(_16043_),
    .S(_16044_));
 FA_X1 _39959_ (.A(_16045_),
    .B(_16046_),
    .CI(_16047_),
    .CO(_16034_),
    .S(_16048_));
 FA_X1 _39960_ (.A(_16021_),
    .B(_16049_),
    .CI(_16043_),
    .CO(_16050_),
    .S(_16051_));
 FA_X1 _39961_ (.A(_16052_),
    .B(_16053_),
    .CI(_16054_),
    .CO(_16055_),
    .S(_16056_));
 FA_X1 _39962_ (.A(net239),
    .B(_16057_),
    .CI(_16058_),
    .CO(_16059_),
    .S(_16060_));
 FA_X1 _39963_ (.A(_16048_),
    .B(_16061_),
    .CI(_16062_),
    .CO(_16063_),
    .S(_16064_));
 FA_X1 _39964_ (.A(_16028_),
    .B(_16065_),
    .CI(_16066_),
    .CO(_16035_),
    .S(_16067_));
 FA_X1 _39965_ (.A(_16068_),
    .B(_16069_),
    .CI(_16070_),
    .CO(_16061_),
    .S(_16071_));
 FA_X1 _39966_ (.A(net44),
    .B(_16072_),
    .CI(_16073_),
    .CO(_16074_),
    .S(_16075_));
 FA_X1 _39967_ (.A(_16076_),
    .B(_16077_),
    .CI(_16044_),
    .CO(_16078_),
    .S(_16079_));
 FA_X1 _39968_ (.A(_16080_),
    .B(_16081_),
    .CI(_16082_),
    .CO(_16083_),
    .S(_16084_));
 FA_X1 _39969_ (.A(_15870_),
    .B(_16085_),
    .CI(_16086_),
    .CO(_16070_),
    .S(_16087_));
 FA_X1 _39970_ (.A(_16071_),
    .B(_16088_),
    .CI(_16089_),
    .CO(_16090_),
    .S(_16091_));
 FA_X1 _39971_ (.A(_16092_),
    .B(_16093_),
    .CI(_16094_),
    .CO(_16062_),
    .S(_16095_));
 FA_X1 _39972_ (.A(_16096_),
    .B(_16097_),
    .CI(_16098_),
    .CO(_16088_),
    .S(_16099_));
 FA_X1 _39973_ (.A(_16100_),
    .B(_16101_),
    .CI(_16102_),
    .CO(_16096_),
    .S(_16103_));
 FA_X1 _39974_ (.A(_16104_),
    .B(_16105_),
    .CI(_16106_),
    .CO(_16107_),
    .S(_16108_));
 FA_X1 _39975_ (.A(net238),
    .B(_16109_),
    .CI(_16110_),
    .CO(_16111_),
    .S(_16112_));
 FA_X1 _39976_ (.A(_16099_),
    .B(_16113_),
    .CI(_16114_),
    .CO(_16115_),
    .S(_16116_));
 FA_X1 _39977_ (.A(_16117_),
    .B(_16118_),
    .CI(_16087_),
    .CO(_16089_),
    .S(_16119_));
 FA_X1 _39978_ (.A(_16120_),
    .B(_16121_),
    .CI(_16122_),
    .CO(_16113_),
    .S(_16123_));
 FA_X1 _39979_ (.A(_16124_),
    .B(_16125_),
    .CI(_16126_),
    .CO(_16127_),
    .S(_16128_));
 FA_X1 _39980_ (.A(_16129_),
    .B(_16130_),
    .CI(_16131_),
    .CO(_16120_),
    .S(_16132_));
 FA_X1 _39981_ (.A(_16133_),
    .B(_16134_),
    .CI(_16135_),
    .CO(_16136_),
    .S(_16137_));
 FA_X1 _39982_ (.A(_16138_),
    .B(_16123_),
    .CI(_16139_),
    .CO(_16140_),
    .S(_16141_));
 FA_X1 _39983_ (.A(_16103_),
    .B(_16142_),
    .CI(_16143_),
    .CO(_16114_),
    .S(_16144_));
 FA_X1 _39984_ (.A(_16145_),
    .B(_16146_),
    .CI(_16147_),
    .CO(_16148_),
    .S(_16149_));
 FA_X1 _39985_ (.A(_16150_),
    .B(_16151_),
    .CI(_16152_),
    .CO(_16146_),
    .S(_16153_));
 FA_X1 _39986_ (.A(_16154_),
    .B(_16155_),
    .CI(_16156_),
    .CO(_16145_),
    .S(_16157_));
 FA_X1 _39987_ (.A(_16158_),
    .B(_16159_),
    .CI(_16160_),
    .CO(_16161_),
    .S(_16162_));
 FA_X1 _39988_ (.A(_16163_),
    .B(_16132_),
    .CI(_16164_),
    .CO(_16139_),
    .S(_16165_));
 FA_X1 _39989_ (.A(_16166_),
    .B(_16167_),
    .CI(_16168_),
    .CO(_16159_),
    .S(_16169_));
 FA_X1 _39990_ (.A(_16170_),
    .B(_16171_),
    .CI(_16172_),
    .CO(_16173_),
    .S(_16174_));
 FA_X1 _39991_ (.A(_16175_),
    .B(_16169_),
    .CI(_16176_),
    .CO(_16177_),
    .S(_16178_));
 FA_X1 _39992_ (.A(_16179_),
    .B(_16180_),
    .CI(_16181_),
    .CO(_16160_),
    .S(_16182_));
 FA_X1 _39993_ (.A(_16183_),
    .B(_16184_),
    .CI(_16185_),
    .CO(_16186_),
    .S(_16187_));
 FA_X1 _39994_ (.A(_16188_),
    .B(_16189_),
    .CI(_16190_),
    .CO(_16191_),
    .S(_16192_));
 FA_X1 _39995_ (.A(_16193_),
    .B(_16194_),
    .CI(_16174_),
    .CO(_16195_),
    .S(_16196_));
 FA_X1 _39996_ (.A(_16197_),
    .B(_16198_),
    .CI(_16199_),
    .CO(_16200_),
    .S(_16201_));
 FA_X1 _39997_ (.A(_16202_),
    .B(_16201_),
    .CI(_16203_),
    .CO(_16204_),
    .S(_16205_));
 FA_X1 _39998_ (.A(_16206_),
    .B(_16207_),
    .CI(_16208_),
    .CO(_16190_),
    .S(_16209_));
 FA_X1 _39999_ (.A(_16210_),
    .B(_16211_),
    .CI(_16212_),
    .CO(_16202_),
    .S(_16213_));
 FA_X1 _40000_ (.A(_16214_),
    .B(_16215_),
    .CI(_16216_),
    .CO(_16217_),
    .S(_16218_));
 FA_X1 _40001_ (.A(_16219_),
    .B(_16220_),
    .CI(_16221_),
    .CO(_16222_),
    .S(_16223_));
 FA_X1 _40002_ (.A(_16224_),
    .B(_16225_),
    .CI(_16226_),
    .CO(_16227_),
    .S(_16228_));
 FA_X1 _40003_ (.A(_16229_),
    .B(_16230_),
    .CI(_16231_),
    .CO(_16232_),
    .S(_16233_));
 FA_X1 _40004_ (.A(_16234_),
    .B(_16235_),
    .CI(_16236_),
    .CO(_16237_),
    .S(_16238_));
 FA_X1 _40005_ (.A(_16239_),
    .B(_16240_),
    .CI(_16241_),
    .CO(_16242_),
    .S(_16243_));
 FA_X1 _40006_ (.A(_16244_),
    .B(_16245_),
    .CI(_16246_),
    .CO(_16247_),
    .S(_16248_));
 FA_X1 _40007_ (.A(_16232_),
    .B(_16248_),
    .CI(_16249_),
    .CO(_16250_),
    .S(_16251_));
 FA_X1 _40008_ (.A(_16252_),
    .B(_16253_),
    .CI(_16254_),
    .CO(_16255_),
    .S(_16256_));
 FA_X1 _40009_ (.A(_16257_),
    .B(_16258_),
    .CI(_16256_),
    .CO(_16259_),
    .S(_16260_));
 FA_X1 _40010_ (.A(_16261_),
    .B(_16262_),
    .CI(_16263_),
    .CO(_16264_),
    .S(_16265_));
 FA_X1 _40011_ (.A(_16266_),
    .B(_16267_),
    .CI(_16242_),
    .CO(_16268_),
    .S(_16269_));
 FA_X1 _40012_ (.A(_16270_),
    .B(_16271_),
    .CI(_16272_),
    .CO(_16273_),
    .S(_16274_));
 FA_X1 _40013_ (.A(_16275_),
    .B(_16276_),
    .CI(_16277_),
    .CO(_16278_),
    .S(_16279_));
 FA_X1 _40014_ (.A(_16280_),
    .B(_16281_),
    .CI(_16282_),
    .CO(_16283_),
    .S(_16284_));
 FA_X1 _40015_ (.A(_16285_),
    .B(_16286_),
    .CI(_16287_),
    .CO(_16288_),
    .S(_16289_));
 FA_X1 _40016_ (.A(_16290_),
    .B(_16289_),
    .CI(_16291_),
    .CO(_16292_),
    .S(_16293_));
 FA_X1 _40017_ (.A(_16294_),
    .B(_16295_),
    .CI(_16296_),
    .CO(_16297_),
    .S(_16298_));
 FA_X1 _40018_ (.A(_16299_),
    .B(_16300_),
    .CI(_16301_),
    .CO(_16302_),
    .S(_16303_));
 FA_X1 _40019_ (.A(_16304_),
    .B(_16305_),
    .CI(_16306_),
    .CO(_16307_),
    .S(_16308_));
 FA_X1 _40020_ (.A(_16298_),
    .B(_16309_),
    .CI(_16310_),
    .CO(_16311_),
    .S(_16312_));
 FA_X1 _40021_ (.A(_16313_),
    .B(_16314_),
    .CI(_16315_),
    .CO(_16316_),
    .S(_16317_));
 FA_X1 _40022_ (.A(_16288_),
    .B(_16317_),
    .CI(_16283_),
    .CO(_16318_),
    .S(_16319_));
 FA_X1 _40023_ (.A(_16320_),
    .B(_16321_),
    .CI(_16322_),
    .CO(_16323_),
    .S(_16324_));
 FA_X1 _40024_ (.A(net92),
    .B(_16325_),
    .CI(_16326_),
    .CO(_16327_),
    .S(_16328_));
 FA_X1 _40025_ (.A(_16329_),
    .B(_16330_),
    .CI(_16328_),
    .CO(_16331_),
    .S(_16332_));
 FA_X1 _40026_ (.A(net232),
    .B(_16333_),
    .CI(_16334_),
    .CO(_16335_),
    .S(_16336_));
 FA_X1 _40027_ (.A(_16337_),
    .B(_16338_),
    .CI(_16339_),
    .CO(_16340_),
    .S(_16341_));
 FA_X1 _40028_ (.A(_16342_),
    .B(_16343_),
    .CI(_16297_),
    .CO(_16344_),
    .S(_16345_));
 FA_X1 _40029_ (.A(_16345_),
    .B(_16316_),
    .CI(_16311_),
    .CO(_16346_),
    .S(_16347_));
 FA_X1 _40030_ (.A(_16348_),
    .B(_16349_),
    .CI(_16350_),
    .CO(_16351_),
    .S(_16352_));
 FA_X1 _40031_ (.A(net93),
    .B(_16353_),
    .CI(_16354_),
    .CO(_16355_),
    .S(_16356_));
 FA_X1 _40032_ (.A(_16357_),
    .B(_16358_),
    .CI(_16359_),
    .CO(_16360_),
    .S(_16361_));
 FA_X1 _40033_ (.A(_15313_),
    .B(_16362_),
    .CI(_16363_),
    .CO(_16364_),
    .S(_16365_));
 FA_X1 _40034_ (.A(_16366_),
    .B(_16361_),
    .CI(_16365_),
    .CO(_16367_),
    .S(_16368_));
 FA_X1 _40035_ (.A(_16369_),
    .B(_16370_),
    .CI(_16371_),
    .CO(_16372_),
    .S(_16373_));
 FA_X1 _40036_ (.A(_16373_),
    .B(_16344_),
    .CI(_16340_),
    .CO(_16374_),
    .S(_16375_));
 FA_X1 _40037_ (.A(_16376_),
    .B(_16377_),
    .CI(_16378_),
    .CO(_16379_),
    .S(_16380_));
 FA_X1 _40038_ (.A(net94),
    .B(_16381_),
    .CI(_16382_),
    .CO(_16383_),
    .S(_16384_));
 FA_X1 _40039_ (.A(_16385_),
    .B(_16384_),
    .CI(_16355_),
    .CO(_16386_),
    .S(_16387_));
 FA_X1 _40040_ (.A(net248),
    .B(_16388_),
    .CI(_16389_),
    .CO(_16390_),
    .S(_16391_));
 FA_X1 _40041_ (.A(_16392_),
    .B(_16393_),
    .CI(_16394_),
    .CO(_16395_),
    .S(_16396_));
 FA_X1 _40042_ (.A(_16397_),
    .B(_16360_),
    .CI(_16364_),
    .CO(_16398_),
    .S(_16399_));
 FA_X1 _40043_ (.A(_16367_),
    .B(_16399_),
    .CI(_16372_),
    .CO(_16400_),
    .S(_16401_));
 FA_X1 _40044_ (.A(_16402_),
    .B(_16403_),
    .CI(_16404_),
    .CO(_16405_),
    .S(_16406_));
 FA_X1 _40045_ (.A(_16398_),
    .B(_16406_),
    .CI(_16395_),
    .CO(_16407_),
    .S(_16408_));
 FA_X1 _40046_ (.A(_15238_),
    .B(_16409_),
    .CI(_16410_),
    .CO(_16411_),
    .S(_16412_));
 FA_X1 _40047_ (.A(net95),
    .B(_16413_),
    .CI(_16414_),
    .CO(_16415_),
    .S(_16416_));
 FA_X1 _40048_ (.A(_16417_),
    .B(_16418_),
    .CI(_16419_),
    .CO(_16420_),
    .S(_16421_));
 FA_X1 _40049_ (.A(_16412_),
    .B(_16422_),
    .CI(_16423_),
    .CO(_16424_),
    .S(_16425_));
 FA_X1 _40050_ (.A(net262),
    .B(_16420_),
    .CI(_16415_),
    .CO(_16426_),
    .S(_16427_));
 FA_X1 _40051_ (.A(_16405_),
    .B(_16428_),
    .CI(_16424_),
    .CO(_16429_),
    .S(_16430_));
 FA_X1 _40052_ (.A(_16431_),
    .B(_16432_),
    .CI(_16433_),
    .CO(_16434_),
    .S(_16435_));
 FA_X1 _40053_ (.A(net96),
    .B(_16436_),
    .CI(_16437_),
    .CO(_16438_),
    .S(_16439_));
 FA_X1 _40054_ (.A(_16440_),
    .B(_16411_),
    .CI(_16441_),
    .CO(_16442_),
    .S(_16443_));
 FA_X1 _40055_ (.A(net270),
    .B(_16444_),
    .CI(_16445_),
    .CO(_16446_),
    .S(_16447_));
 FA_X1 _40056_ (.A(_16448_),
    .B(_16449_),
    .CI(_16442_),
    .CO(_16450_),
    .S(_16451_));
 FA_X1 _40057_ (.A(net97),
    .B(_16452_),
    .CI(_16453_),
    .CO(_16454_),
    .S(_16455_));
 FA_X1 _40058_ (.A(_16456_),
    .B(_16457_),
    .CI(_16458_),
    .CO(_16459_),
    .S(_16460_));
 FA_X1 _40059_ (.A(_15196_),
    .B(_16461_),
    .CI(_16462_),
    .CO(_16463_),
    .S(_16464_));
 FA_X1 _40060_ (.A(net98),
    .B(_16465_),
    .CI(_16466_),
    .CO(_16467_),
    .S(_16468_));
 FA_X1 _40061_ (.A(_16469_),
    .B(_16459_),
    .CI(_16470_),
    .CO(_16471_),
    .S(_16472_));
 FA_X1 _40062_ (.A(_15651_),
    .B(_16473_),
    .CI(_16474_),
    .CO(_16475_),
    .S(_16476_));
 FA_X1 _40063_ (.A(net67),
    .B(_16477_),
    .CI(_16478_),
    .CO(_16479_),
    .S(_16480_));
 FA_X1 _40064_ (.A(_16481_),
    .B(_15761_),
    .CI(_16482_),
    .CO(_16483_),
    .S(_16484_));
 FA_X1 _40065_ (.A(_16485_),
    .B(_16486_),
    .CI(_16487_),
    .CO(_16488_),
    .S(_16489_));
 FA_X1 _40066_ (.A(net274),
    .B(_16467_),
    .CI(_16490_),
    .CO(_16491_),
    .S(_16492_));
 FA_X1 _40067_ (.A(net101),
    .B(net275),
    .CI(_16493_),
    .CO(_16494_),
    .S(_16495_));
 FA_X1 _40068_ (.A(net53),
    .B(net243),
    .CI(_16496_),
    .CO(_16497_),
    .S(_16498_));
 FA_X1 _40069_ (.A(net242),
    .B(_16499_),
    .CI(_16500_),
    .CO(_16501_),
    .S(_16502_));
 FA_X1 _40070_ (.A(net52),
    .B(_16503_),
    .CI(_16504_),
    .CO(_16505_),
    .S(_16506_));
 FA_X1 _40071_ (.A(net51),
    .B(_16507_),
    .CI(_16508_),
    .CO(_16500_),
    .S(_16509_));
 FA_X1 _40072_ (.A(_16510_),
    .B(_16511_),
    .CI(_16012_),
    .CO(_16512_),
    .S(_16513_));
 FA_X1 _40073_ (.A(_15964_),
    .B(_16514_),
    .CI(_16515_),
    .CO(_16516_),
    .S(_16517_));
 FA_X1 _40074_ (.A(_16518_),
    .B(_16519_),
    .CI(_16520_),
    .CO(_16521_),
    .S(_16522_));
 FA_X1 _40075_ (.A(_16523_),
    .B(_16524_),
    .CI(_16525_),
    .CO(_16526_),
    .S(_16527_));
 FA_X1 _40076_ (.A(_16528_),
    .B(_16529_),
    .CI(_16530_),
    .CO(_16531_),
    .S(_16532_));
 FA_X1 _40077_ (.A(_16533_),
    .B(_16534_),
    .CI(_16535_),
    .CO(_16536_),
    .S(_16537_));
 FA_X1 _40078_ (.A(_16538_),
    .B(_16539_),
    .CI(_16540_),
    .CO(_16541_),
    .S(_16542_));
 FA_X1 _40079_ (.A(_16543_),
    .B(_16542_),
    .CI(_16544_),
    .CO(_16545_),
    .S(_16546_));
 FA_X1 _40080_ (.A(_16547_),
    .B(_16548_),
    .CI(_16549_),
    .CO(_16523_),
    .S(_16550_));
 FA_X1 _40081_ (.A(_16551_),
    .B(_16552_),
    .CI(_16553_),
    .CO(_16544_),
    .S(_16554_));
 FA_X1 _40082_ (.A(_16555_),
    .B(_16556_),
    .CI(_16557_),
    .CO(_16558_),
    .S(_16559_));
 FA_X1 _40083_ (.A(_16560_),
    .B(_16561_),
    .CI(_16562_),
    .CO(_16563_),
    .S(_16564_));
 FA_X1 _40084_ (.A(net221),
    .B(net275),
    .CI(_16565_),
    .CO(_16566_),
    .S(_16567_));
 FA_X1 _40085_ (.A(net160),
    .B(_16568_),
    .CI(_16569_),
    .CO(_16570_),
    .S(_16571_));
 FA_X1 _40086_ (.A(_16572_),
    .B(_16573_),
    .CI(_16574_),
    .CO(_16575_),
    .S(_16576_));
 FA_X1 _40087_ (.A(net100),
    .B(_16577_),
    .CI(_16578_),
    .CO(_16579_),
    .S(_16580_));
 FA_X1 _40088_ (.A(_16581_),
    .B(_16582_),
    .CI(_16583_),
    .CO(_16584_),
    .S(_16585_));
 FA_X1 _40089_ (.A(_16571_),
    .B(_16579_),
    .CI(_16586_),
    .CO(_16587_),
    .S(_16588_));
 FA_X1 _40090_ (.A(net248),
    .B(_16589_),
    .CI(_16590_),
    .CO(_16591_),
    .S(_16592_));
 FA_X1 _40091_ (.A(_16576_),
    .B(_16593_),
    .CI(_16594_),
    .CO(_16595_),
    .S(_16596_));
 FA_X1 _40092_ (.A(net171),
    .B(_16597_),
    .CI(_16598_),
    .CO(_16599_),
    .S(_16600_));
 FA_X1 _40093_ (.A(_15238_),
    .B(_16601_),
    .CI(_16602_),
    .CO(_16603_),
    .S(_16604_));
 FA_X1 _40094_ (.A(_16605_),
    .B(_16606_),
    .CI(_16607_),
    .CO(_16608_),
    .S(_16609_));
 FA_X1 _40095_ (.A(_16610_),
    .B(_16604_),
    .CI(_16611_),
    .CO(_16612_),
    .S(_16613_));
 FA_X1 _40096_ (.A(_16614_),
    .B(_16615_),
    .CI(_16616_),
    .CO(_16593_),
    .S(_16617_));
 FA_X1 _40097_ (.A(net1),
    .B(_16618_),
    .CI(_16619_),
    .CO(_16620_),
    .S(_16621_));
 FA_X1 _40098_ (.A(_16622_),
    .B(_16623_),
    .CI(_16624_),
    .CO(_16625_),
    .S(_16626_));
 FA_X1 _40099_ (.A(_16627_),
    .B(_16628_),
    .CI(_16629_),
    .CO(_16615_),
    .S(_16630_));
 FA_X1 _40100_ (.A(_15313_),
    .B(_16631_),
    .CI(_16632_),
    .CO(_16616_),
    .S(_16633_));
 FA_X1 _40101_ (.A(_16634_),
    .B(_16635_),
    .CI(_16636_),
    .CO(_16637_),
    .S(_16638_));
 FA_X1 _40102_ (.A(_16639_),
    .B(_16640_),
    .CI(_16641_),
    .CO(_16635_),
    .S(_16642_));
 FA_X1 _40103_ (.A(_16643_),
    .B(_16644_),
    .CI(_16645_),
    .CO(_16636_),
    .S(_16646_));
 FA_X1 _40104_ (.A(_16647_),
    .B(_16648_),
    .CI(_16649_),
    .CO(_16650_),
    .S(_16651_));
 FA_X1 _40105_ (.A(_16652_),
    .B(_16653_),
    .CI(_16654_),
    .CO(_16655_),
    .S(_16656_));
 FA_X1 _40106_ (.A(_16657_),
    .B(_16658_),
    .CI(_16659_),
    .CO(_16660_),
    .S(_16661_));
 FA_X1 _40107_ (.A(_16662_),
    .B(_16663_),
    .CI(_16664_),
    .CO(_16665_),
    .S(_16666_));
 FA_X1 _40108_ (.A(_16667_),
    .B(_16656_),
    .CI(_16668_),
    .CO(_16669_),
    .S(_16670_));
 FA_X1 _40109_ (.A(_16671_),
    .B(_16672_),
    .CI(_16673_),
    .CO(_16647_),
    .S(_16674_));
 FA_X1 _40110_ (.A(_16675_),
    .B(_16676_),
    .CI(_16677_),
    .CO(_16678_),
    .S(_16679_));
 FA_X1 _40111_ (.A(_16680_),
    .B(_16681_),
    .CI(_16682_),
    .CO(_16683_),
    .S(_16684_));
 FA_X1 _40112_ (.A(_16685_),
    .B(_16686_),
    .CI(_16687_),
    .CO(_16688_),
    .S(_16689_));
 FA_X1 _40113_ (.A(_14689_),
    .B(_16690_),
    .CI(_16691_),
    .CO(_16692_),
    .S(_16693_));
 FA_X1 _40114_ (.A(_16694_),
    .B(_14655_),
    .CI(_16695_),
    .CO(_14661_),
    .S(_16696_));
 FA_X1 _40115_ (.A(_16697_),
    .B(_16698_),
    .CI(_16699_),
    .CO(_16700_),
    .S(_16701_));
 FA_X1 _40116_ (.A(_16702_),
    .B(_16703_),
    .CI(_16704_),
    .CO(_16697_),
    .S(_16705_));
 FA_X1 _40117_ (.A(_16706_),
    .B(_16707_),
    .CI(_16708_),
    .CO(_16699_),
    .S(_16709_));
 FA_X1 _40118_ (.A(_16710_),
    .B(_16711_),
    .CI(_16712_),
    .CO(_16713_),
    .S(_16714_));
 FA_X1 _40119_ (.A(_16715_),
    .B(_14698_),
    .CI(_16716_),
    .CO(_16691_),
    .S(_16717_));
 FA_X1 _40120_ (.A(_16718_),
    .B(_16719_),
    .CI(_16720_),
    .CO(_16712_),
    .S(_16721_));
 FA_X1 _40121_ (.A(_16722_),
    .B(_16723_),
    .CI(_16724_),
    .CO(_16725_),
    .S(_16726_));
 FA_X1 _40122_ (.A(net254),
    .B(_16727_),
    .CI(_16479_),
    .CO(_16728_),
    .S(_16729_));
 FA_X1 _40123_ (.A(_16721_),
    .B(_16536_),
    .CI(_16730_),
    .CO(_16731_),
    .S(_16732_));
 FA_X1 _40124_ (.A(_16733_),
    .B(_16734_),
    .CI(_16735_),
    .CO(_16711_),
    .S(_16736_));
 FA_X1 _40125_ (.A(net219),
    .B(_16737_),
    .CI(_16738_),
    .CO(_16739_),
    .S(_16740_));
 FA_X1 _40126_ (.A(net242),
    .B(_16741_),
    .CI(_16742_),
    .CO(_16743_),
    .S(_16744_));
 FA_X1 _40127_ (.A(net218),
    .B(_16746_),
    .CI(_16747_),
    .CO(_16742_),
    .S(_16748_));
 FA_X1 _40128_ (.A(net217),
    .B(_16749_),
    .CI(_16750_),
    .CO(_16751_),
    .S(_16752_));
 FA_X1 _40129_ (.A(net213),
    .B(_16753_),
    .CI(_16754_),
    .CO(_16755_),
    .S(_16756_));
 FA_X1 _40130_ (.A(net214),
    .B(_16757_),
    .CI(_16758_),
    .CO(_16759_),
    .S(_16760_));
 FA_X1 _40131_ (.A(_16761_),
    .B(_16762_),
    .CI(_16763_),
    .CO(_16764_),
    .S(_16765_));
 FA_X1 _40132_ (.A(_16760_),
    .B(_16755_),
    .CI(_16766_),
    .CO(_16767_),
    .S(_16768_));
 FA_X1 _40133_ (.A(_16769_),
    .B(_16770_),
    .CI(_16771_),
    .CO(_16772_),
    .S(_16773_));
 FA_X1 _40134_ (.A(net239),
    .B(_16774_),
    .CI(_16775_),
    .CO(_16776_),
    .S(_16777_));
 FA_X1 _40135_ (.A(_16778_),
    .B(_16765_),
    .CI(_16779_),
    .CO(_16780_),
    .S(_16781_));
 FA_X1 _40136_ (.A(net215),
    .B(_16782_),
    .CI(_16783_),
    .CO(_16784_),
    .S(_16785_));
 FA_X1 _40137_ (.A(_15915_),
    .B(_16786_),
    .CI(_16787_),
    .CO(_16788_),
    .S(_16789_));
 FA_X1 _40138_ (.A(_16790_),
    .B(_16791_),
    .CI(_16792_),
    .CO(_16793_),
    .S(_16794_));
 FA_X1 _40139_ (.A(_16789_),
    .B(_16795_),
    .CI(_16796_),
    .CO(_16797_),
    .S(_16798_));
 FA_X1 _40140_ (.A(_16799_),
    .B(_16800_),
    .CI(_16801_),
    .CO(_16778_),
    .S(_16802_));
 FA_X1 _40141_ (.A(net212),
    .B(_16803_),
    .CI(_16804_),
    .CO(_16805_),
    .S(_16806_));
 FA_X1 _40142_ (.A(_16807_),
    .B(_16808_),
    .CI(_16809_),
    .CO(_16810_),
    .S(_16811_));
 FA_X1 _40143_ (.A(_16756_),
    .B(_16812_),
    .CI(_16813_),
    .CO(_16814_),
    .S(_16815_));
 FA_X1 _40144_ (.A(_15870_),
    .B(_16816_),
    .CI(_16817_),
    .CO(_16801_),
    .S(_16818_));
 FA_X1 _40145_ (.A(_16819_),
    .B(_16820_),
    .CI(_16821_),
    .CO(_16822_),
    .S(_16823_));
 FA_X1 _40146_ (.A(_16824_),
    .B(_16825_),
    .CI(_16826_),
    .CO(_16827_),
    .S(_16828_));
 FA_X1 _40147_ (.A(_16829_),
    .B(_16830_),
    .CI(_16823_),
    .CO(_16831_),
    .S(_16832_));
 FA_X1 _40148_ (.A(_16833_),
    .B(_16834_),
    .CI(_16835_),
    .CO(_16836_),
    .S(_16837_));
 FA_X1 _40149_ (.A(_16838_),
    .B(_16839_),
    .CI(_16840_),
    .CO(_16841_),
    .S(_16842_));
 FA_X1 _40150_ (.A(_16843_),
    .B(_16844_),
    .CI(_16845_),
    .CO(_16846_),
    .S(_16847_));
 FA_X1 _40151_ (.A(_16848_),
    .B(_16849_),
    .CI(_16850_),
    .CO(_16851_),
    .S(_16852_));
 FA_X1 _40152_ (.A(net270),
    .B(_16853_),
    .CI(_16854_),
    .CO(_16855_),
    .S(_16856_));
 FA_X1 _40153_ (.A(_16857_),
    .B(_16858_),
    .CI(_16859_),
    .CO(_16860_),
    .S(_16861_));
 FA_X1 _40154_ (.A(net199),
    .B(_16862_),
    .CI(_16863_),
    .CO(_16864_),
    .S(_16865_));
 FA_X1 _40155_ (.A(_16866_),
    .B(_16867_),
    .CI(_16868_),
    .CO(_16869_),
    .S(_16870_));
 FA_X1 _40156_ (.A(net200),
    .B(_16871_),
    .CI(_16872_),
    .CO(_16873_),
    .S(_16874_));
 FA_X1 _40157_ (.A(_16875_),
    .B(_16876_),
    .CI(_16877_),
    .CO(_16878_),
    .S(_16879_));
 FA_X1 _40158_ (.A(net262),
    .B(_16880_),
    .CI(_16881_),
    .CO(_16882_),
    .S(_16883_));
 FA_X1 _40159_ (.A(net197),
    .B(_16884_),
    .CI(_16885_),
    .CO(_16886_),
    .S(_16887_));
 FA_X1 _40160_ (.A(_15238_),
    .B(_16888_),
    .CI(_16889_),
    .CO(_16890_),
    .S(_16891_));
 FA_X1 _40161_ (.A(net198),
    .B(_16892_),
    .CI(_16893_),
    .CO(_16881_),
    .S(_16894_));
 FA_X1 _40162_ (.A(_16895_),
    .B(_16896_),
    .CI(_16897_),
    .CO(_16880_),
    .S(_16898_));
 FA_X1 _40163_ (.A(_16899_),
    .B(_16900_),
    .CI(_16901_),
    .CO(_16902_),
    .S(_16903_));
 FA_X1 _40164_ (.A(_16904_),
    .B(_16905_),
    .CI(_16906_),
    .CO(_16900_),
    .S(_16907_));
 FA_X1 _40165_ (.A(_16908_),
    .B(_16909_),
    .CI(_16910_),
    .CO(_16911_),
    .S(_16912_));
 FA_X1 _40166_ (.A(_16913_),
    .B(_16914_),
    .CI(_16915_),
    .CO(_16916_),
    .S(_16917_));
 FA_X1 _40167_ (.A(_16903_),
    .B(_16918_),
    .CI(_16919_),
    .CO(_16920_),
    .S(_16921_));
 FA_X1 _40168_ (.A(_16922_),
    .B(_16923_),
    .CI(_16924_),
    .CO(_16925_),
    .S(_16926_));
 FA_X1 _40169_ (.A(net195),
    .B(_16927_),
    .CI(_16928_),
    .CO(_16929_),
    .S(_16930_));
 FA_X1 _40170_ (.A(_16931_),
    .B(_16932_),
    .CI(_16930_),
    .CO(_16933_),
    .S(_16934_));
 FA_X1 _40171_ (.A(net232),
    .B(_16935_),
    .CI(_16936_),
    .CO(_16937_),
    .S(_16938_));
 FA_X1 _40172_ (.A(_16939_),
    .B(_16940_),
    .CI(_16941_),
    .CO(_16942_),
    .S(_16943_));
 FA_X1 _40173_ (.A(_16944_),
    .B(_16945_),
    .CI(_16946_),
    .CO(_16947_),
    .S(_16948_));
 FA_X1 _40174_ (.A(_16949_),
    .B(_16950_),
    .CI(_16951_),
    .CO(_16944_),
    .S(_16952_));
 FA_X1 _40175_ (.A(_16953_),
    .B(_16954_),
    .CI(_16955_),
    .CO(_16946_),
    .S(_16956_));
 FA_X1 _40176_ (.A(_16957_),
    .B(_16958_),
    .CI(_16959_),
    .CO(_16960_),
    .S(_16961_));
 FA_X1 _40177_ (.A(_16962_),
    .B(_16961_),
    .CI(_16963_),
    .CO(_16964_),
    .S(_16965_));
 FA_X1 _40178_ (.A(_16966_),
    .B(_16967_),
    .CI(_16968_),
    .CO(_16969_),
    .S(_16970_));
 FA_X1 _40179_ (.A(_16971_),
    .B(_16972_),
    .CI(_16973_),
    .CO(_16962_),
    .S(_16974_));
 FA_X1 _40180_ (.A(_16975_),
    .B(_16976_),
    .CI(_16977_),
    .CO(_16978_),
    .S(_16979_));
 FA_X1 _40181_ (.A(net266),
    .B(_16980_),
    .CI(_16981_),
    .CO(_16982_),
    .S(_16983_));
 FA_X1 _40182_ (.A(net186),
    .B(_16985_),
    .CI(_16986_),
    .CO(_16981_),
    .S(_16987_));
 FA_X1 _40183_ (.A(net185),
    .B(_16988_),
    .CI(_16989_),
    .CO(_16990_),
    .S(_16991_));
 FA_X1 _40184_ (.A(net180),
    .B(_16992_),
    .CI(_16993_),
    .CO(_16994_),
    .S(_16995_));
 FA_X1 _40185_ (.A(net182),
    .B(_16996_),
    .CI(_16997_),
    .CO(_16998_),
    .S(_16999_));
 FA_X1 _40186_ (.A(_17000_),
    .B(_17001_),
    .CI(_17002_),
    .CO(_17003_),
    .S(_17004_));
 FA_X1 _40187_ (.A(_16999_),
    .B(_16994_),
    .CI(_17005_),
    .CO(_17006_),
    .S(_17007_));
 FA_X1 _40188_ (.A(_17008_),
    .B(_17009_),
    .CI(_17010_),
    .CO(_17011_),
    .S(_17012_));
 FA_X1 _40189_ (.A(net263),
    .B(_17013_),
    .CI(_17014_),
    .CO(_17015_),
    .S(_17016_));
 FA_X1 _40190_ (.A(_17017_),
    .B(_17004_),
    .CI(_17018_),
    .CO(_17019_),
    .S(_17020_));
 FA_X1 _40191_ (.A(net183),
    .B(_17021_),
    .CI(_17022_),
    .CO(_17023_),
    .S(_17024_));
 FA_X1 _40192_ (.A(_14888_),
    .B(_17025_),
    .CI(_17026_),
    .CO(_17027_),
    .S(_17028_));
 FA_X1 _40193_ (.A(_17029_),
    .B(_17030_),
    .CI(_17031_),
    .CO(_17032_),
    .S(_17033_));
 FA_X1 _40194_ (.A(_17034_),
    .B(_17028_),
    .CI(_17035_),
    .CO(_17036_),
    .S(_17037_));
 FA_X1 _40195_ (.A(net179),
    .B(_17038_),
    .CI(_17039_),
    .CO(_17040_),
    .S(_17041_));
 FA_X1 _40196_ (.A(_17042_),
    .B(_17043_),
    .CI(_17044_),
    .CO(_17017_),
    .S(_17045_));
 FA_X1 _40197_ (.A(_17046_),
    .B(_17047_),
    .CI(_16995_),
    .CO(_17048_),
    .S(_17049_));
 FA_X1 _40198_ (.A(_17050_),
    .B(_17051_),
    .CI(_17052_),
    .CO(_17053_),
    .S(_17054_));
 FA_X1 _40199_ (.A(_14841_),
    .B(_17055_),
    .CI(_17056_),
    .CO(_17044_),
    .S(_17057_));
 FA_X1 _40200_ (.A(_17058_),
    .B(_17059_),
    .CI(_17060_),
    .CO(_17061_),
    .S(_17062_));
 FA_X1 _40201_ (.A(_17063_),
    .B(_17064_),
    .CI(_17065_),
    .CO(_17066_),
    .S(_17067_));
 FA_X1 _40202_ (.A(_17068_),
    .B(_17069_),
    .CI(_17070_),
    .CO(_17071_),
    .S(_17072_));
 FA_X1 _40203_ (.A(_17073_),
    .B(_17067_),
    .CI(_17074_),
    .CO(_17075_),
    .S(_17076_));
 FA_X1 _40204_ (.A(_17077_),
    .B(_17078_),
    .CI(_17079_),
    .CO(_17080_),
    .S(_17081_));
 FA_X1 _40205_ (.A(_17082_),
    .B(_17083_),
    .CI(_17084_),
    .CO(_17077_),
    .S(_17085_));
 FA_X1 _40206_ (.A(_17086_),
    .B(_17087_),
    .CI(_17088_),
    .CO(_17079_),
    .S(_17089_));
 FA_X1 _40207_ (.A(_17090_),
    .B(_17091_),
    .CI(_17092_),
    .CO(_17093_),
    .S(_17094_));
 FA_X1 _40208_ (.A(_17095_),
    .B(_17096_),
    .CI(_17097_),
    .CO(_17091_),
    .S(_17098_));
 FA_X1 _40209_ (.A(_17099_),
    .B(_17100_),
    .CI(_17101_),
    .CO(_17102_),
    .S(_17103_));
 FA_X1 _40210_ (.A(_17104_),
    .B(_17105_),
    .CI(_17106_),
    .CO(_17107_),
    .S(_17108_));
 FA_X1 _40211_ (.A(_17109_),
    .B(_17110_),
    .CI(_17111_),
    .CO(_17112_),
    .S(_17113_));
 FA_X1 _40212_ (.A(net254),
    .B(_17114_),
    .CI(_17115_),
    .CO(_17116_),
    .S(_17117_));
 FA_X1 _40213_ (.A(net170),
    .B(_17118_),
    .CI(_17119_),
    .CO(_17120_),
    .S(_17121_));
 FA_X1 _40214_ (.A(net169),
    .B(_17122_),
    .CI(_17123_),
    .CO(_17115_),
    .S(_17124_));
 FA_X1 _40215_ (.A(net168),
    .B(_17125_),
    .CI(_17126_),
    .CO(_17127_),
    .S(_17128_));
 FA_X1 _40216_ (.A(_15412_),
    .B(_17129_),
    .CI(_17130_),
    .CO(_17131_),
    .S(_17132_));
 FA_X1 _40217_ (.A(net166),
    .B(_17133_),
    .CI(_17134_),
    .CO(_17135_),
    .S(_17136_));
 FA_X1 _40218_ (.A(_17137_),
    .B(_17138_),
    .CI(_17139_),
    .CO(_17140_),
    .S(_17141_));
 FA_X1 _40219_ (.A(_17142_),
    .B(_17132_),
    .CI(_17143_),
    .CO(_17144_),
    .S(_17145_));
 FA_X1 _40220_ (.A(net165),
    .B(_17146_),
    .CI(_17147_),
    .CO(_17148_),
    .S(_17149_));
 FA_X1 _40221_ (.A(_17150_),
    .B(_17151_),
    .CI(_17152_),
    .CO(_17153_),
    .S(_17154_));
 FA_X1 _40222_ (.A(net164),
    .B(_17155_),
    .CI(_17156_),
    .CO(_17157_),
    .S(_17158_));
 FA_X1 _40223_ (.A(_17159_),
    .B(_17160_),
    .CI(_17161_),
    .CO(_17162_),
    .S(_17163_));
 FA_X1 _40224_ (.A(_17149_),
    .B(_17157_),
    .CI(_17164_),
    .CO(_17165_),
    .S(_17166_));
 FA_X1 _40225_ (.A(net251),
    .B(_17167_),
    .CI(_17168_),
    .CO(_17169_),
    .S(_17170_));
 FA_X1 _40226_ (.A(_17154_),
    .B(_17171_),
    .CI(_17172_),
    .CO(_17173_),
    .S(_17174_));
 FA_X1 _40227_ (.A(net163),
    .B(_17175_),
    .CI(_17176_),
    .CO(_17177_),
    .S(_17178_));
 FA_X1 _40228_ (.A(_17179_),
    .B(_17180_),
    .CI(_17181_),
    .CO(_17171_),
    .S(_17182_));
 FA_X1 _40229_ (.A(_17183_),
    .B(_17184_),
    .CI(_17185_),
    .CO(_17186_),
    .S(_17187_));
 FA_X1 _40230_ (.A(_17188_),
    .B(_17189_),
    .CI(_17190_),
    .CO(_17180_),
    .S(_17191_));
 FA_X1 _40231_ (.A(_14677_),
    .B(_17192_),
    .CI(_17193_),
    .CO(_17181_),
    .S(_17194_));
 FA_X1 _40232_ (.A(_17195_),
    .B(_17196_),
    .CI(_17197_),
    .CO(_17198_),
    .S(_17199_));
 FA_X1 _40233_ (.A(_17200_),
    .B(_17201_),
    .CI(_17202_),
    .CO(_17203_),
    .S(_17204_));
 FA_X1 _40234_ (.A(_17205_),
    .B(_17206_),
    .CI(_17207_),
    .CO(_17208_),
    .S(_17209_));
 FA_X1 _40235_ (.A(_17204_),
    .B(_17210_),
    .CI(_17211_),
    .CO(_17212_),
    .S(_17213_));
 FA_X1 _40236_ (.A(_17214_),
    .B(_17215_),
    .CI(_17216_),
    .CO(_17217_),
    .S(_17218_));
 FA_X1 _40237_ (.A(_17219_),
    .B(_17220_),
    .CI(_17221_),
    .CO(_17222_),
    .S(_17223_));
 FA_X1 _40238_ (.A(_17224_),
    .B(_17225_),
    .CI(_17226_),
    .CO(_17227_),
    .S(_17228_));
 FA_X1 _40239_ (.A(_17218_),
    .B(_17229_),
    .CI(_17230_),
    .CO(_17231_),
    .S(_17232_));
 FA_X1 _40240_ (.A(_17233_),
    .B(_17234_),
    .CI(_17235_),
    .CO(_17229_),
    .S(_17236_));
 FA_X1 _40241_ (.A(_17237_),
    .B(_17238_),
    .CI(_17239_),
    .CO(_17240_),
    .S(_17241_));
 FA_X1 _40242_ (.A(_17242_),
    .B(_17243_),
    .CI(_17244_),
    .CO(_17245_),
    .S(_17246_));
 FA_X1 _40243_ (.A(_17247_),
    .B(_17248_),
    .CI(_17249_),
    .CO(_17250_),
    .S(_17251_));
 FA_X1 _40244_ (.A(_17252_),
    .B(_17253_),
    .CI(_17254_),
    .CO(_17255_),
    .S(_17256_));
 FA_X1 _40245_ (.A(_17257_),
    .B(_17258_),
    .CI(_17259_),
    .CO(_17252_),
    .S(_17260_));
 FA_X1 _40246_ (.A(_17261_),
    .B(_17262_),
    .CI(_17263_),
    .CO(_17254_),
    .S(_17264_));
 FA_X1 _40247_ (.A(_17265_),
    .B(_17266_),
    .CI(_17267_),
    .CO(_17268_),
    .S(_17269_));
 FA_X1 _40248_ (.A(_17270_),
    .B(_17271_),
    .CI(_17272_),
    .CO(_17273_),
    .S(_17274_));
 FA_X1 _40249_ (.A(_17275_),
    .B(_17276_),
    .CI(_17277_),
    .CO(_17278_),
    .S(_17279_));
 FA_X1 _40250_ (.A(_17280_),
    .B(_17281_),
    .CI(_17282_),
    .CO(_17283_),
    .S(_17284_));
 FA_X1 _40251_ (.A(_17285_),
    .B(_17279_),
    .CI(_17286_),
    .CO(_17287_),
    .S(_17288_));
 FA_X1 _40252_ (.A(_17289_),
    .B(_17290_),
    .CI(_17291_),
    .CO(_17266_),
    .S(_17292_));
 FA_X1 _40253_ (.A(_17293_),
    .B(_17294_),
    .CI(_17295_),
    .CO(_17296_),
    .S(_17297_));
 FA_X1 _40254_ (.A(net69),
    .B(_17298_),
    .CI(_17299_),
    .CO(_17300_),
    .S(_17301_));
 FA_X1 _40255_ (.A(_17302_),
    .B(_17303_),
    .CI(_17304_),
    .CO(_17305_),
    .S(_17306_));
 FA_X1 _40256_ (.A(_17307_),
    .B(_17308_),
    .CI(_17309_),
    .CO(_17303_),
    .S(_17310_));
 FA_X1 _40257_ (.A(_17311_),
    .B(_17312_),
    .CI(_17313_),
    .CO(_17314_),
    .S(_17315_));
 FA_X1 _40258_ (.A(net238),
    .B(_17316_),
    .CI(_17317_),
    .CO(_17318_),
    .S(_17319_));
 FA_X1 _40259_ (.A(_17306_),
    .B(_17320_),
    .CI(_17321_),
    .CO(_17322_),
    .S(_17323_));
 FA_X1 _40260_ (.A(net80),
    .B(_17324_),
    .CI(_17325_),
    .CO(_17326_),
    .S(_17327_));
 FA_X1 _40261_ (.A(_17327_),
    .B(_17328_),
    .CI(_17329_),
    .CO(_17330_),
    .S(_17331_));
 FA_X1 _40262_ (.A(_17332_),
    .B(_17333_),
    .CI(_17334_),
    .CO(_17335_),
    .S(_17336_));
 FA_X1 _40263_ (.A(_15870_),
    .B(_17337_),
    .CI(_17338_),
    .CO(_17339_),
    .S(_17340_));
 FA_X1 _40264_ (.A(_17341_),
    .B(_17342_),
    .CI(_17340_),
    .CO(_17343_),
    .S(_17344_));
 FA_X1 _40265_ (.A(_17278_),
    .B(_17345_),
    .CI(_17346_),
    .CO(_17320_),
    .S(_17347_));
 FA_X1 _40266_ (.A(_17348_),
    .B(_17349_),
    .CI(_17350_),
    .CO(_17351_),
    .S(_17352_));
 FA_X1 _40267_ (.A(net242),
    .B(_17353_),
    .CI(_17354_),
    .CO(_17355_),
    .S(_17356_));
 FA_X1 _40268_ (.A(net131),
    .B(_17358_),
    .CI(_17359_),
    .CO(_17354_),
    .S(_17360_));
 FA_X1 _40269_ (.A(net120),
    .B(_17361_),
    .CI(_17362_),
    .CO(_17363_),
    .S(_17364_));
 FA_X1 _40270_ (.A(_17365_),
    .B(_17366_),
    .CI(_17367_),
    .CO(_17368_),
    .S(_17369_));
 FA_X1 _40271_ (.A(_17370_),
    .B(_17371_),
    .CI(_17372_),
    .CO(_17373_),
    .S(_17374_));
 FA_X1 _40272_ (.A(_17375_),
    .B(_17376_),
    .CI(_17297_),
    .CO(_17377_),
    .S(_17378_));
 FA_X1 _40273_ (.A(_17379_),
    .B(_17380_),
    .CI(_17381_),
    .CO(_17382_),
    .S(_17383_));
 FA_X1 _40274_ (.A(_17384_),
    .B(_17385_),
    .CI(_17386_),
    .CO(_17387_),
    .S(_17388_));
 FA_X1 _40275_ (.A(net241),
    .B(_17389_),
    .CI(_17390_),
    .CO(_17391_),
    .S(_17392_));
 FA_X1 _40276_ (.A(_17393_),
    .B(_17394_),
    .CI(_17395_),
    .CO(_17396_),
    .S(_17397_));
 FA_X1 _40277_ (.A(net110),
    .B(_17398_),
    .CI(_17399_),
    .CO(_17400_),
    .S(_17401_));
 FA_X1 _40278_ (.A(_17402_),
    .B(_17403_),
    .CI(_17404_),
    .CO(_17405_),
    .S(_17406_));
 FA_X1 _40279_ (.A(net240),
    .B(_17407_),
    .CI(_17408_),
    .CO(_17409_),
    .S(_17410_));
 FA_X1 _40280_ (.A(net89),
    .B(_17411_),
    .CI(_17412_),
    .CO(_17413_),
    .S(_17414_));
 FA_X1 _40281_ (.A(net99),
    .B(_17415_),
    .CI(_17416_),
    .CO(_17408_),
    .S(_17417_));
 FA_X1 _40282_ (.A(_15915_),
    .B(_17418_),
    .CI(_17419_),
    .CO(_17420_),
    .S(_17421_));
 FA_X1 _40283_ (.A(_17422_),
    .B(_17423_),
    .CI(_17424_),
    .CO(_17407_),
    .S(_17425_));
 FA_X1 _40284_ (.A(_17426_),
    .B(_17427_),
    .CI(_17428_),
    .CO(_17429_),
    .S(_17430_));
 FA_X1 _40285_ (.A(_17431_),
    .B(_17432_),
    .CI(_17433_),
    .CO(_17434_),
    .S(_17435_));
 FA_X1 _40286_ (.A(_17436_),
    .B(_17437_),
    .CI(_17438_),
    .CO(_17439_),
    .S(_17440_));
 FA_X1 _40287_ (.A(net229),
    .B(_17441_),
    .CI(_17442_),
    .CO(_17443_),
    .S(_17444_));
 FA_X1 _40288_ (.A(_17445_),
    .B(_17446_),
    .CI(_17447_),
    .CO(_17448_),
    .S(_17449_));
 FA_X1 _40289_ (.A(net228),
    .B(_17450_),
    .CI(_17451_),
    .CO(_17452_),
    .S(_17453_));
 FA_X1 _40290_ (.A(_17454_),
    .B(_17455_),
    .CI(_17456_),
    .CO(_17457_),
    .S(_17458_));
 FA_X1 _40291_ (.A(_17459_),
    .B(_17460_),
    .CI(_17444_),
    .CO(_17461_),
    .S(_17462_));
 FA_X1 _40292_ (.A(_14677_),
    .B(_17463_),
    .CI(_17464_),
    .CO(_17447_),
    .S(_17465_));
 FA_X1 _40293_ (.A(_17449_),
    .B(_17466_),
    .CI(_17467_),
    .CO(_17468_),
    .S(_17469_));
 FA_X1 _40294_ (.A(_17470_),
    .B(_17471_),
    .CI(_17472_),
    .CO(_17473_),
    .S(_17474_));
 FA_X1 _40295_ (.A(net230),
    .B(_17475_),
    .CI(_17476_),
    .CO(_17477_),
    .S(_17478_));
 FA_X1 _40296_ (.A(_17479_),
    .B(_17443_),
    .CI(_17478_),
    .CO(_17480_),
    .S(_17481_));
 FA_X1 _40297_ (.A(net251),
    .B(_17482_),
    .CI(_17483_),
    .CO(_17484_),
    .S(_17485_));
 FA_X1 _40298_ (.A(_17486_),
    .B(_17487_),
    .CI(_17488_),
    .CO(_17489_),
    .S(_17490_));
 FA_X1 _40299_ (.A(_17491_),
    .B(_17492_),
    .CI(_17493_),
    .CO(_17466_),
    .S(_17494_));
 FA_X1 _40300_ (.A(_17495_),
    .B(_17496_),
    .CI(_17497_),
    .CO(_17498_),
    .S(_17499_));
 FA_X1 _40301_ (.A(_17500_),
    .B(_17501_),
    .CI(_17502_),
    .CO(_17492_),
    .S(_17503_));
 FA_X1 _40302_ (.A(net250),
    .B(_17504_),
    .CI(_17505_),
    .CO(_17506_),
    .S(_17507_));
 FA_X1 _40303_ (.A(_17508_),
    .B(_17509_),
    .CI(_17510_),
    .CO(_17511_),
    .S(_17512_));
 FA_X1 _40304_ (.A(_17513_),
    .B(_17514_),
    .CI(_17515_),
    .CO(_17508_),
    .S(_17516_));
 FA_X1 _40305_ (.A(_17517_),
    .B(_17518_),
    .CI(_17519_),
    .CO(_17520_),
    .S(_17521_));
 FA_X1 _40306_ (.A(net238),
    .B(_17522_),
    .CI(_17523_),
    .CO(_17524_),
    .S(_17525_));
 FA_X1 _40307_ (.A(_17526_),
    .B(_17512_),
    .CI(_17527_),
    .CO(_17528_),
    .S(_17529_));
 FA_X1 _40308_ (.A(_17530_),
    .B(_17531_),
    .CI(_16818_),
    .CO(_17532_),
    .S(_17533_));
 FA_X1 _40309_ (.A(_17534_),
    .B(_17535_),
    .CI(_17536_),
    .CO(_17526_),
    .S(_17537_));
 FA_X1 _40310_ (.A(_17538_),
    .B(_17539_),
    .CI(_17540_),
    .CO(_17541_),
    .S(_17542_));
 FA_X1 _40311_ (.A(_17543_),
    .B(_17544_),
    .CI(_17545_),
    .CO(_17534_),
    .S(_17546_));
 FA_X1 _40312_ (.A(_17547_),
    .B(_17548_),
    .CI(_17549_),
    .CO(_17550_),
    .S(_17551_));
 FA_X1 _40313_ (.A(_17552_),
    .B(_17553_),
    .CI(_17554_),
    .CO(_17555_),
    .S(_17556_));
 FA_X1 _40314_ (.A(_17557_),
    .B(_17558_),
    .CI(_17559_),
    .CO(_17560_),
    .S(_17561_));
 FA_X1 _40315_ (.A(_17556_),
    .B(_17562_),
    .CI(_17563_),
    .CO(_17564_),
    .S(_17565_));
 FA_X1 _40316_ (.A(_17566_),
    .B(_17567_),
    .CI(_17568_),
    .CO(_17569_),
    .S(_17570_));
 FA_X1 _40317_ (.A(_17571_),
    .B(_17572_),
    .CI(_17573_),
    .CO(_17574_),
    .S(_17575_));
 FA_X1 _40318_ (.A(_17576_),
    .B(_17577_),
    .CI(_17057_),
    .CO(_17578_),
    .S(_17579_));
 FA_X1 _40319_ (.A(_17580_),
    .B(_17581_),
    .CI(_17582_),
    .CO(_17583_),
    .S(_17584_));
 FA_X1 _40320_ (.A(_17585_),
    .B(_17586_),
    .CI(_17041_),
    .CO(_17587_),
    .S(_17588_));
 FA_X1 _40321_ (.A(_17589_),
    .B(_17590_),
    .CI(_17591_),
    .CO(_17592_),
    .S(_17593_));
 FA_X1 _40322_ (.A(net261),
    .B(_17594_),
    .CI(_17595_),
    .CO(_17596_),
    .S(_17597_));
 FA_X1 _40323_ (.A(_17584_),
    .B(_17598_),
    .CI(_17599_),
    .CO(_17600_),
    .S(_17601_));
 FA_X1 _40324_ (.A(_17066_),
    .B(_17602_),
    .CI(_17603_),
    .CO(_17598_),
    .S(_17604_));
 FA_X1 _40325_ (.A(net253),
    .B(_17605_),
    .CI(_17606_),
    .CO(_17607_),
    .S(_17608_));
 FA_X1 _40326_ (.A(_17609_),
    .B(_17610_),
    .CI(_17611_),
    .CO(_17612_),
    .S(_17613_));
 FA_X1 _40327_ (.A(net167),
    .B(_17614_),
    .CI(_17615_),
    .CO(_17616_),
    .S(_17617_));
 FA_X1 _40328_ (.A(_17618_),
    .B(_17619_),
    .CI(_17620_),
    .CO(_17621_),
    .S(_17622_));
 FA_X1 _40329_ (.A(_17623_),
    .B(_17624_),
    .CI(_17625_),
    .CO(_17626_),
    .S(_17627_));
 FA_X1 _40330_ (.A(net252),
    .B(_17140_),
    .CI(_17135_),
    .CO(_17628_),
    .S(_17629_));
 FA_X1 _40331_ (.A(_17630_),
    .B(_17631_),
    .CI(_17632_),
    .CO(_17633_),
    .S(_17634_));
 FA_X1 _40332_ (.A(_17635_),
    .B(_17636_),
    .CI(_17637_),
    .CO(_17638_),
    .S(_17639_));
 FA_X1 _40333_ (.A(net201),
    .B(_17640_),
    .CI(_17641_),
    .CO(_17642_),
    .S(_17643_));
 FA_X1 _40334_ (.A(net190),
    .B(_17644_),
    .CI(_17645_),
    .CO(_17646_),
    .S(_17647_));
 FA_X1 _40335_ (.A(_17648_),
    .B(_17649_),
    .CI(_17650_),
    .CO(_17651_),
    .S(_17652_));
 FA_X1 _40336_ (.A(_15196_),
    .B(_17653_),
    .CI(_17654_),
    .CO(_17655_),
    .S(_17656_));
 FA_X1 _40337_ (.A(net270),
    .B(_17657_),
    .CI(_17658_),
    .CO(_17659_),
    .S(_17660_));
 FA_X1 _40338_ (.A(_17661_),
    .B(_17662_),
    .CI(_17663_),
    .CO(_17664_),
    .S(_17665_));
 FA_X1 _40339_ (.A(net181),
    .B(_17666_),
    .CI(_17667_),
    .CO(_17668_),
    .S(_17669_));
 FA_X1 _40340_ (.A(_17670_),
    .B(_17671_),
    .CI(_17672_),
    .CO(_17673_),
    .S(_17674_));
 FA_X1 _40341_ (.A(net266),
    .B(_17675_),
    .CI(_17676_),
    .CO(_17677_),
    .S(_17678_));
 FA_X1 _40342_ (.A(net19),
    .B(_17680_),
    .CI(_17681_),
    .CO(_17675_),
    .S(_17682_));
 FA_X1 _40343_ (.A(net18),
    .B(_17683_),
    .CI(_17684_),
    .CO(_17685_),
    .S(_17686_));
 FA_X1 _40344_ (.A(net16),
    .B(_17687_),
    .CI(_17688_),
    .CO(_17689_),
    .S(_17690_));
 FA_X1 _40345_ (.A(_14888_),
    .B(_17691_),
    .CI(_17692_),
    .CO(_17693_),
    .S(_17694_));
 FA_X1 _40346_ (.A(_17695_),
    .B(_17696_),
    .CI(_17697_),
    .CO(_17698_),
    .S(_17699_));
 FA_X1 _40347_ (.A(_17694_),
    .B(_17700_),
    .CI(_17701_),
    .CO(_17702_),
    .S(_17703_));
 FA_X1 _40348_ (.A(net14),
    .B(_17704_),
    .CI(_17705_),
    .CO(_17706_),
    .S(_17707_));
 FA_X1 _40349_ (.A(net15),
    .B(_17708_),
    .CI(_17709_),
    .CO(_17710_),
    .S(_17711_));
 FA_X1 _40350_ (.A(_17712_),
    .B(_17713_),
    .CI(_17714_),
    .CO(_17715_),
    .S(_17716_));
 FA_X1 _40351_ (.A(_17717_),
    .B(_17706_),
    .CI(_17711_),
    .CO(_17718_),
    .S(_17719_));
 FA_X1 _40352_ (.A(_17720_),
    .B(_17721_),
    .CI(_17722_),
    .CO(_17723_),
    .S(_17724_));
 FA_X1 _40353_ (.A(net263),
    .B(_17725_),
    .CI(_17726_),
    .CO(_17727_),
    .S(_17728_));
 FA_X1 _40354_ (.A(_17729_),
    .B(_17730_),
    .CI(_17716_),
    .CO(_17731_),
    .S(_17732_));
 FA_X1 _40355_ (.A(_17733_),
    .B(_17734_),
    .CI(_17735_),
    .CO(_17729_),
    .S(_17736_));
 FA_X1 _40356_ (.A(net13),
    .B(_17737_),
    .CI(_17738_),
    .CO(_17739_),
    .S(_17740_));
 FA_X1 _40357_ (.A(_17741_),
    .B(_17742_),
    .CI(_17707_),
    .CO(_17743_),
    .S(_17744_));
 FA_X1 _40358_ (.A(_17745_),
    .B(_17746_),
    .CI(_17747_),
    .CO(_17748_),
    .S(_17749_));
 FA_X1 _40359_ (.A(_14841_),
    .B(_17750_),
    .CI(_17751_),
    .CO(_17735_),
    .S(_17752_));
 FA_X1 _40360_ (.A(_17753_),
    .B(_17754_),
    .CI(_17752_),
    .CO(_17755_),
    .S(_17756_));
 FA_X1 _40361_ (.A(_17757_),
    .B(_17758_),
    .CI(_17759_),
    .CO(_17760_),
    .S(_17761_));
 FA_X1 _40362_ (.A(_17762_),
    .B(_17763_),
    .CI(_17740_),
    .CO(_17764_),
    .S(_17765_));
 FA_X1 _40363_ (.A(_17766_),
    .B(_17767_),
    .CI(_17768_),
    .CO(_17769_),
    .S(_17770_));
 FA_X1 _40364_ (.A(net261),
    .B(_17771_),
    .CI(_17772_),
    .CO(_17773_),
    .S(_17774_));
 FA_X1 _40365_ (.A(_17761_),
    .B(_17775_),
    .CI(_17776_),
    .CO(_17777_),
    .S(_17778_));
 FA_X1 _40366_ (.A(_17779_),
    .B(_17780_),
    .CI(_17781_),
    .CO(_17775_),
    .S(_17782_));
 FA_X1 _40367_ (.A(_17783_),
    .B(_17784_),
    .CI(_17785_),
    .CO(_17786_),
    .S(_17787_));
 FA_X1 _40368_ (.A(_17788_),
    .B(_17789_),
    .CI(_17790_),
    .CO(_17780_),
    .S(_17791_));
 FA_X1 _40369_ (.A(_17792_),
    .B(_17793_),
    .CI(_17794_),
    .CO(_17795_),
    .S(_17796_));
 FA_X1 _40370_ (.A(_17797_),
    .B(_17798_),
    .CI(_17799_),
    .CO(_17800_),
    .S(_17801_));
 FA_X1 _40371_ (.A(_17802_),
    .B(_17803_),
    .CI(_17801_),
    .CO(_17804_),
    .S(_17805_));
 FA_X1 _40372_ (.A(_17806_),
    .B(_17807_),
    .CI(_17808_),
    .CO(_17809_),
    .S(_17810_));
 FA_X1 _40373_ (.A(_17811_),
    .B(_17812_),
    .CI(_17813_),
    .CO(_17814_),
    .S(_17815_));
 FA_X1 _40374_ (.A(_17816_),
    .B(_17817_),
    .CI(_17818_),
    .CO(_17819_),
    .S(_17820_));
 FA_X1 _40375_ (.A(net5),
    .B(net255),
    .CI(_17821_),
    .CO(_17822_),
    .S(_17823_));
 FA_X1 _40376_ (.A(_17824_),
    .B(_17825_),
    .CI(_17826_),
    .CO(_17827_),
    .S(_17828_));
 FA_X1 _40377_ (.A(net2),
    .B(_17829_),
    .CI(_17830_),
    .CO(_17831_),
    .S(_17832_));
 FA_X1 _40378_ (.A(_17833_),
    .B(_17834_),
    .CI(_17835_),
    .CO(_17836_),
    .S(_17837_));
 FA_X1 _40379_ (.A(net252),
    .B(_17838_),
    .CI(_17839_),
    .CO(_17840_),
    .S(_17841_));
 FA_X1 _40380_ (.A(_15412_),
    .B(_17842_),
    .CI(_17843_),
    .CO(_17834_),
    .S(_17844_));
 FA_X1 _40381_ (.A(net231),
    .B(_17845_),
    .CI(_17846_),
    .CO(_17839_),
    .S(_17847_));
 FA_X1 _40382_ (.A(_17848_),
    .B(_17849_),
    .CI(_17850_),
    .CO(_17838_),
    .S(_17851_));
 FA_X1 _40383_ (.A(_17852_),
    .B(_17853_),
    .CI(_17854_),
    .CO(_17855_),
    .S(_17856_));
 FA_X1 _40384_ (.A(_17857_),
    .B(_17858_),
    .CI(_17859_),
    .CO(_17853_),
    .S(_17860_));
 FA_X1 _40385_ (.A(_17861_),
    .B(_17862_),
    .CI(_17863_),
    .CO(_17864_),
    .S(_17865_));
 FA_X1 _40386_ (.A(_17866_),
    .B(_17867_),
    .CI(_17868_),
    .CO(_17862_),
    .S(_17869_));
 FA_X1 _40387_ (.A(_17870_),
    .B(_17871_),
    .CI(_17872_),
    .CO(_17873_),
    .S(_17874_));
 FA_X1 _40388_ (.A(_17875_),
    .B(_17876_),
    .CI(_17877_),
    .CO(_17878_),
    .S(_17879_));
 FA_X1 _40389_ (.A(_17865_),
    .B(_17880_),
    .CI(_17881_),
    .CO(_17882_),
    .S(_17883_));
 FA_X1 _40390_ (.A(_17884_),
    .B(_17503_),
    .CI(_17885_),
    .CO(_17886_),
    .S(_17887_));
 FA_X1 _40391_ (.A(_17888_),
    .B(_17889_),
    .CI(_17890_),
    .CO(_17891_),
    .S(_17892_));
 FA_X1 _40392_ (.A(_17893_),
    .B(_17894_),
    .CI(_17895_),
    .CO(_17889_),
    .S(_17896_));
 FA_X1 _40393_ (.A(_17897_),
    .B(_17898_),
    .CI(_17899_),
    .CO(_17890_),
    .S(_17900_));
 FA_X1 _40394_ (.A(_17901_),
    .B(_17902_),
    .CI(_17903_),
    .CO(_17904_),
    .S(_17905_));
 FA_X1 _40395_ (.A(_17906_),
    .B(_17907_),
    .CI(_17908_),
    .CO(_17909_),
    .S(_17910_));
 FA_X1 _40396_ (.A(_17905_),
    .B(_17911_),
    .CI(_17912_),
    .CO(_17913_),
    .S(_17914_));
 FA_X1 _40397_ (.A(_17915_),
    .B(_17916_),
    .CI(_17917_),
    .CO(_17918_),
    .S(_17919_));
 FA_X1 _40398_ (.A(_17920_),
    .B(_17921_),
    .CI(_17922_),
    .CO(_17923_),
    .S(_17924_));
 FA_X1 _40399_ (.A(_17925_),
    .B(_17926_),
    .CI(_17927_),
    .CO(_17928_),
    .S(_17929_));
 FA_X1 _40400_ (.A(_17930_),
    .B(_17931_),
    .CI(_17932_),
    .CO(_17933_),
    .S(_17934_));
 FA_X1 _40401_ (.A(_17935_),
    .B(_17936_),
    .CI(_17937_),
    .CO(_17926_),
    .S(_17938_));
 FA_X1 _40402_ (.A(net232),
    .B(_17939_),
    .CI(_17940_),
    .CO(_17941_),
    .S(_17942_));
 FA_X1 _40403_ (.A(_17943_),
    .B(_17929_),
    .CI(_17944_),
    .CO(_17945_),
    .S(_17946_));
 FA_X1 _40404_ (.A(_16633_),
    .B(_16630_),
    .CI(_17947_),
    .CO(_17948_),
    .S(_17949_));
 FA_X1 _40405_ (.A(_16655_),
    .B(_17950_),
    .CI(_17951_),
    .CO(_17944_),
    .S(_17952_));
 FA_X1 _40406_ (.A(_17953_),
    .B(_17954_),
    .CI(_17955_),
    .CO(_17956_),
    .S(_17957_));
 FA_X1 _40407_ (.A(_17326_),
    .B(_17414_),
    .CI(_17958_),
    .CO(_17959_),
    .S(_17960_));
 FA_X1 _40408_ (.A(_17961_),
    .B(_17962_),
    .CI(_17963_),
    .CO(_17964_),
    .S(_17965_));
 FA_X1 _40409_ (.A(net239),
    .B(_17966_),
    .CI(_17967_),
    .CO(_17968_),
    .S(_17969_));
 FA_X1 _40410_ (.A(_17957_),
    .B(_17970_),
    .CI(_17971_),
    .CO(_17972_),
    .S(_17973_));
 FA_X1 _40411_ (.A(_17974_),
    .B(_17421_),
    .CI(_17975_),
    .CO(_17976_),
    .S(_17977_));
 FA_X1 _40412_ (.A(_17978_),
    .B(_17339_),
    .CI(_17979_),
    .CO(_17970_),
    .S(_17980_));
 FA_X1 _40413_ (.A(_17241_),
    .B(_17981_),
    .CI(_17982_),
    .CO(_17983_),
    .S(_17984_));
 FA_X1 _40414_ (.A(_17985_),
    .B(_17986_),
    .CI(_17987_),
    .CO(_17988_),
    .S(_17989_));
 FA_X1 _40415_ (.A(_17990_),
    .B(_17991_),
    .CI(_17992_),
    .CO(_17993_),
    .S(_17994_));
 FA_X1 _40416_ (.A(_17995_),
    .B(_17996_),
    .CI(_17997_),
    .CO(_17998_),
    .S(_17999_));
 FA_X1 _40417_ (.A(_17194_),
    .B(_17191_),
    .CI(_18000_),
    .CO(_18001_),
    .S(_18002_));
 FA_X1 _40418_ (.A(_18003_),
    .B(_18004_),
    .CI(_18005_),
    .CO(_18006_),
    .S(_18007_));
 FA_X1 _40419_ (.A(_18008_),
    .B(_18009_),
    .CI(_18010_),
    .CO(_18011_),
    .S(_18012_));
 FA_X1 _40420_ (.A(_18013_),
    .B(_18014_),
    .CI(_17178_),
    .CO(_18015_),
    .S(_18016_));
 FA_X1 _40421_ (.A(net250),
    .B(_18017_),
    .CI(_18018_),
    .CO(_18019_),
    .S(_18020_));
 FA_X1 _40422_ (.A(_18007_),
    .B(_18021_),
    .CI(_18022_),
    .CO(_18023_),
    .S(_18024_));
 FA_X1 _40423_ (.A(_18025_),
    .B(_17203_),
    .CI(_18026_),
    .CO(_18021_),
    .S(_18027_));
 FA_X1 _40424_ (.A(_18028_),
    .B(_18029_),
    .CI(_17103_),
    .CO(_18030_),
    .S(_18031_));
 FA_X1 _40425_ (.A(_18032_),
    .B(_18033_),
    .CI(_18034_),
    .CO(_18035_),
    .S(_18036_));
 FA_X1 _40426_ (.A(_18037_),
    .B(_18038_),
    .CI(_18039_),
    .CO(_18040_),
    .S(_18041_));
 FA_X1 _40427_ (.A(_18042_),
    .B(_18043_),
    .CI(_18044_),
    .CO(_18045_),
    .S(_18046_));
 FA_X1 _40428_ (.A(_18047_),
    .B(_18048_),
    .CI(_18049_),
    .CO(_18050_),
    .S(_18051_));
 FA_X1 _40429_ (.A(net265),
    .B(_18052_),
    .CI(_18053_),
    .CO(_18054_),
    .S(_18055_));
 FA_X1 _40430_ (.A(_18056_),
    .B(_18057_),
    .CI(_18058_),
    .CO(_18059_),
    .S(_18060_));
 FA_X1 _40431_ (.A(net184),
    .B(_18061_),
    .CI(_18062_),
    .CO(_18063_),
    .S(_18064_));
 FA_X1 _40432_ (.A(_18065_),
    .B(_18066_),
    .CI(_18067_),
    .CO(_18068_),
    .S(_18069_));
 FA_X1 _40433_ (.A(net264),
    .B(_17032_),
    .CI(_17023_),
    .CO(_18070_),
    .S(_18071_));
 FA_X1 _40434_ (.A(_18072_),
    .B(_18073_),
    .CI(_18074_),
    .CO(_18075_),
    .S(_18076_));
 FA_X1 _40435_ (.A(net196),
    .B(_18077_),
    .CI(_18078_),
    .CO(_18079_),
    .S(_18080_));
 FA_X1 _40436_ (.A(_18081_),
    .B(_18082_),
    .CI(_18083_),
    .CO(_18084_),
    .S(_18085_));
 FA_X1 _40437_ (.A(_18086_),
    .B(_18087_),
    .CI(_18088_),
    .CO(_18089_),
    .S(_18090_));
 FA_X1 _40438_ (.A(_16887_),
    .B(_18079_),
    .CI(_18091_),
    .CO(_18092_),
    .S(_18093_));
 FA_X1 _40439_ (.A(net248),
    .B(_18094_),
    .CI(_18095_),
    .CO(_18096_),
    .S(_18097_));
 FA_X1 _40440_ (.A(_18085_),
    .B(_18098_),
    .CI(_18099_),
    .CO(_18100_),
    .S(_18101_));
 FA_X1 _40441_ (.A(_18102_),
    .B(_16891_),
    .CI(_18103_),
    .CO(_18104_),
    .S(_18105_));
 FA_X1 _40442_ (.A(_18106_),
    .B(_18107_),
    .CI(_18108_),
    .CO(_18098_),
    .S(_18109_));
 FA_X1 _40443_ (.A(_18110_),
    .B(_18111_),
    .CI(_18112_),
    .CO(_18113_),
    .S(_18114_));
 FA_X1 _40444_ (.A(_18115_),
    .B(_18116_),
    .CI(_18117_),
    .CO(_18107_),
    .S(_18118_));
 FA_X1 _40445_ (.A(_15313_),
    .B(_18119_),
    .CI(_18120_),
    .CO(_18108_),
    .S(_18121_));
 FA_X1 _40446_ (.A(_18122_),
    .B(_18123_),
    .CI(_18124_),
    .CO(_18125_),
    .S(_18126_));
 FA_X1 _40447_ (.A(_18127_),
    .B(_18128_),
    .CI(_18129_),
    .CO(_18130_),
    .S(_18131_));
 FA_X1 _40448_ (.A(net241),
    .B(_18132_),
    .CI(_18133_),
    .CO(_18134_),
    .S(_18135_));
 FA_X1 _40449_ (.A(_18136_),
    .B(_18137_),
    .CI(_18138_),
    .CO(_18139_),
    .S(_18140_));
 FA_X1 _40450_ (.A(net216),
    .B(_18141_),
    .CI(_18142_),
    .CO(_18143_),
    .S(_18144_));
 FA_X1 _40451_ (.A(_18145_),
    .B(_18146_),
    .CI(_18147_),
    .CO(_18148_),
    .S(_18149_));
 FA_X1 _40452_ (.A(_18150_),
    .B(_18151_),
    .CI(_18152_),
    .CO(_18153_),
    .S(_18154_));
 FA_X1 _40453_ (.A(net240),
    .B(_16793_),
    .CI(_16784_),
    .CO(_18155_),
    .S(_18156_));
 FA_X1 _40454_ (.A(_18157_),
    .B(_18158_),
    .CI(_18159_),
    .CO(_18160_),
    .S(_18161_));
 FA_X1 _40455_ (.A(_18162_),
    .B(_18161_),
    .CI(_18163_),
    .CO(_18164_),
    .S(_18165_));
 FA_X1 _40456_ (.A(_18166_),
    .B(_18167_),
    .CI(_18168_),
    .CO(_18169_),
    .S(_18170_));
 FA_X1 _40457_ (.A(_18171_),
    .B(_18172_),
    .CI(_18173_),
    .CO(_18162_),
    .S(_18174_));
 FA_X1 _40458_ (.A(_15651_),
    .B(_18175_),
    .CI(_18176_),
    .CO(_18177_),
    .S(_18178_));
 FA_X1 _40459_ (.A(net4),
    .B(_18179_),
    .CI(_18180_),
    .CO(_18181_),
    .S(_18182_));
 FA_X1 _40460_ (.A(net3),
    .B(_18183_),
    .CI(_18184_),
    .CO(_18185_),
    .S(_18186_));
 FA_X1 _40461_ (.A(_18187_),
    .B(_18188_),
    .CI(_18189_),
    .CO(_18190_),
    .S(_18191_));
 FA_X1 _40462_ (.A(net253),
    .B(_18192_),
    .CI(_18193_),
    .CO(_18194_),
    .S(_18195_));
 FA_X1 _40463_ (.A(_18196_),
    .B(_17791_),
    .CI(_18197_),
    .CO(_18198_),
    .S(_18199_));
 FA_X1 _40464_ (.A(_18200_),
    .B(_18201_),
    .CI(_18202_),
    .CO(_18203_),
    .S(_18204_));
 FA_X1 _40465_ (.A(_18205_),
    .B(_18206_),
    .CI(_18207_),
    .CO(_18200_),
    .S(_18208_));
 FA_X1 _40466_ (.A(_18209_),
    .B(_18210_),
    .CI(_18211_),
    .CO(_18202_),
    .S(_18212_));
 FA_X1 _40467_ (.A(_18213_),
    .B(_18214_),
    .CI(_18215_),
    .CO(_18216_),
    .S(_18217_));
 FA_X1 _40468_ (.A(_18218_),
    .B(_18219_),
    .CI(_18220_),
    .CO(_18213_),
    .S(_18221_));
 FA_X1 _40469_ (.A(_18222_),
    .B(_18223_),
    .CI(_18224_),
    .CO(_18225_),
    .S(_18226_));
 FA_X1 _40470_ (.A(_18227_),
    .B(_18228_),
    .CI(_18229_),
    .CO(_18230_),
    .S(_18231_));
 FA_X1 _40471_ (.A(_18232_),
    .B(_16679_),
    .CI(_18233_),
    .CO(_18234_),
    .S(_18235_));
 FA_X1 _40472_ (.A(_18236_),
    .B(_18237_),
    .CI(_18238_),
    .CO(_18239_),
    .S(_18240_));
 FA_X1 _40473_ (.A(net274),
    .B(_18241_),
    .CI(_18242_),
    .CO(_18243_),
    .S(_18244_));
 FA_X1 _40474_ (.A(net203),
    .B(_18245_),
    .CI(_18246_),
    .CO(_18247_),
    .S(_18248_));
 FA_X1 _40475_ (.A(net202),
    .B(_18249_),
    .CI(_18250_),
    .CO(_18242_),
    .S(_18251_));
 FA_X1 _40476_ (.A(_18252_),
    .B(_18253_),
    .CI(_18254_),
    .CO(_18255_),
    .S(_18256_));
 FA_X1 _40477_ (.A(net265),
    .B(_18257_),
    .CI(_18258_),
    .CO(_18259_),
    .S(_18260_));
 FA_X1 _40478_ (.A(_18261_),
    .B(_18262_),
    .CI(_18263_),
    .CO(_18264_),
    .S(_18265_));
 FA_X1 _40479_ (.A(net17),
    .B(_18266_),
    .CI(_18267_),
    .CO(_18268_),
    .S(_18269_));
 FA_X1 _40480_ (.A(_18270_),
    .B(_18271_),
    .CI(_18272_),
    .CO(_18273_),
    .S(_18274_));
 FA_X1 _40481_ (.A(net264),
    .B(_17698_),
    .CI(_17689_),
    .CO(_18275_),
    .S(_18276_));
 FA_X1 _40482_ (.A(_18277_),
    .B(_18278_),
    .CI(_18279_),
    .CO(_18280_),
    .S(_18281_));
 FA_X1 _40483_ (.A(_18282_),
    .B(_18283_),
    .CI(_18169_),
    .CO(_18284_),
    .S(_18285_));
 FA_X1 _40484_ (.A(_18286_),
    .B(_18287_),
    .CI(_18288_),
    .CO(_17912_),
    .S(_18289_));
 FA_X1 _40485_ (.A(_18290_),
    .B(_17918_),
    .CI(_17904_),
    .CO(_18291_),
    .S(_18292_));
 FA_X1 _40486_ (.A(_18293_),
    .B(_17869_),
    .CI(_18294_),
    .CO(_17880_),
    .S(_18295_));
 FA_X1 _40487_ (.A(_17494_),
    .B(_17864_),
    .CI(_17886_),
    .CO(_18296_),
    .S(_18297_));
 FA_X1 _40488_ (.A(_18298_),
    .B(_18299_),
    .CI(_17465_),
    .CO(_17467_),
    .S(_18300_));
 FA_X1 _40489_ (.A(_17860_),
    .B(_17448_),
    .CI(_17489_),
    .CO(_18301_),
    .S(_18302_));
 FA_X1 _40490_ (.A(_17844_),
    .B(_18303_),
    .CI(_18304_),
    .CO(_17854_),
    .S(_18305_));
 FA_X1 _40491_ (.A(_18306_),
    .B(_18307_),
    .CI(_18308_),
    .CO(_18189_),
    .S(_18309_));
 FA_X1 _40492_ (.A(_18310_),
    .B(_18311_),
    .CI(_17836_),
    .CO(_18312_),
    .S(_18313_));
 FA_X1 _40493_ (.A(_18314_),
    .B(_18315_),
    .CI(_18316_),
    .CO(_18317_),
    .S(_18318_));
 FA_X1 _40494_ (.A(net254),
    .B(_18319_),
    .CI(_18181_),
    .CO(_18320_),
    .S(_18321_));
 FA_X1 _40495_ (.A(_18322_),
    .B(_18323_),
    .CI(_18324_),
    .CO(_18325_),
    .S(_18326_));
 FA_X1 _40496_ (.A(_18327_),
    .B(_18328_),
    .CI(_18329_),
    .CO(_17813_),
    .S(_18330_));
 FA_X1 _40497_ (.A(_18331_),
    .B(_17820_),
    .CI(_17434_),
    .CO(_18332_),
    .S(_18333_));
 FA_X1 _40498_ (.A(_18334_),
    .B(_18335_),
    .CI(_18336_),
    .CO(_18215_),
    .S(_18337_));
 FA_X1 _40499_ (.A(_18338_),
    .B(_18221_),
    .CI(_18339_),
    .CO(_18340_),
    .S(_18341_));
 FA_X1 _40500_ (.A(_18342_),
    .B(_18343_),
    .CI(_18344_),
    .CO(_17776_),
    .S(_18345_));
 FA_X1 _40501_ (.A(_17782_),
    .B(_18346_),
    .CI(_18198_),
    .CO(_18347_),
    .S(_18348_));
 FA_X1 _40502_ (.A(_18349_),
    .B(_18350_),
    .CI(_18351_),
    .CO(_17730_),
    .S(_18352_));
 FA_X1 _40503_ (.A(_17736_),
    .B(_17760_),
    .CI(_17755_),
    .CO(_18353_),
    .S(_18354_));
 FA_X1 _40504_ (.A(_18355_),
    .B(_18356_),
    .CI(_17693_),
    .CO(_18272_),
    .S(_18357_));
 FA_X1 _40505_ (.A(_18358_),
    .B(_17715_),
    .CI(_17702_),
    .CO(_18359_),
    .S(_18360_));
 FA_X1 _40506_ (.A(_14944_),
    .B(_18361_),
    .CI(_18362_),
    .CO(_17679_),
    .S(_18363_));
 FA_X1 _40507_ (.A(_18364_),
    .B(_18365_),
    .CI(_18255_),
    .CO(_18366_),
    .S(_18367_));
 FA_X1 _40508_ (.A(net21),
    .B(net267),
    .CI(_18368_),
    .CO(_18369_),
    .S(_18370_));
 FA_X1 _40509_ (.A(_18371_),
    .B(_18372_),
    .CI(_18373_),
    .CO(_18374_),
    .S(_18375_));
 FA_X1 _40510_ (.A(_18376_),
    .B(_18377_),
    .CI(_16969_),
    .CO(_18378_),
    .S(_18379_));
 FA_X1 _40511_ (.A(_18380_),
    .B(_18381_),
    .CI(_17561_),
    .CO(_18382_),
    .S(_18383_));
 FA_X1 _40512_ (.A(_18384_),
    .B(_17555_),
    .CI(_17569_),
    .CO(_18385_),
    .S(_18386_));
 FA_X1 _40513_ (.A(_18387_),
    .B(_16907_),
    .CI(_18388_),
    .CO(_16919_),
    .S(_18389_));
 FA_X1 _40514_ (.A(_18390_),
    .B(_18391_),
    .CI(_18392_),
    .CO(_18393_),
    .S(_18394_));
 FA_X1 _40515_ (.A(_16902_),
    .B(_18394_),
    .CI(_16942_),
    .CO(_18395_),
    .S(_18396_));
 FA_X1 _40516_ (.A(_18121_),
    .B(_18118_),
    .CI(_18397_),
    .CO(_18398_),
    .S(_18399_));
 FA_X1 _40517_ (.A(_18109_),
    .B(_18393_),
    .CI(_18398_),
    .CO(_18400_),
    .S(_18401_));
 FA_X1 _40518_ (.A(_18402_),
    .B(_18403_),
    .CI(_18404_),
    .CO(_18099_),
    .S(_18405_));
 FA_X1 _40519_ (.A(_16890_),
    .B(_18406_),
    .CI(_18407_),
    .CO(_16868_),
    .S(_18408_));
 FA_X1 _40520_ (.A(_18409_),
    .B(_18084_),
    .CI(_18104_),
    .CO(_18410_),
    .S(_18411_));
 FA_X1 _40521_ (.A(_18412_),
    .B(_16878_),
    .CI(_18413_),
    .CO(_18414_),
    .S(_18415_));
 FA_X1 _40522_ (.A(_15196_),
    .B(_18416_),
    .CI(_18417_),
    .CO(_18418_),
    .S(_18419_));
 FA_X1 _40523_ (.A(net204),
    .B(net275),
    .CI(_18420_),
    .CO(_18421_),
    .S(_18422_));
 FA_X1 _40524_ (.A(_18423_),
    .B(_18424_),
    .CI(_18425_),
    .CO(_18426_),
    .S(_18427_));
 FA_X1 _40525_ (.A(_18428_),
    .B(_18429_),
    .CI(_18430_),
    .CO(_18431_),
    .S(_18432_));
 FA_X1 _40526_ (.A(_18125_),
    .B(_18432_),
    .CI(_18433_),
    .CO(_18434_),
    .S(_18435_));
 FA_X1 _40527_ (.A(_18436_),
    .B(_18437_),
    .CI(_18438_),
    .CO(_18439_),
    .S(_18440_));
 FA_X1 _40528_ (.A(_18441_),
    .B(_18442_),
    .CI(_18439_),
    .CO(_18443_),
    .S(_18444_));
 FA_X1 _40529_ (.A(_18445_),
    .B(_18446_),
    .CI(_18447_),
    .CO(_16830_),
    .S(_18448_));
 FA_X1 _40530_ (.A(_16836_),
    .B(_18449_),
    .CI(_16841_),
    .CO(_18450_),
    .S(_18451_));
 FA_X1 _40531_ (.A(_16846_),
    .B(_18452_),
    .CI(_16822_),
    .CO(_18453_),
    .S(_18454_));
 FA_X1 _40532_ (.A(_17546_),
    .B(_18455_),
    .CI(_18456_),
    .CO(_18457_),
    .S(_18458_));
 FA_X1 _40533_ (.A(_17537_),
    .B(_18459_),
    .CI(_18457_),
    .CO(_18460_),
    .S(_18461_));
 FA_X1 _40534_ (.A(_17516_),
    .B(_18462_),
    .CI(_18463_),
    .CO(_17527_),
    .S(_18464_));
 FA_X1 _40535_ (.A(_16802_),
    .B(_17511_),
    .CI(_17532_),
    .CO(_18465_),
    .S(_18466_));
 FA_X1 _40536_ (.A(_18467_),
    .B(_18468_),
    .CI(_18469_),
    .CO(_16779_),
    .S(_18470_));
 FA_X1 _40537_ (.A(_16764_),
    .B(_18471_),
    .CI(_16797_),
    .CO(_18472_),
    .S(_18473_));
 FA_X1 _40538_ (.A(_16788_),
    .B(_18474_),
    .CI(_18475_),
    .CO(_18147_),
    .S(_18476_));
 FA_X1 _40539_ (.A(_18477_),
    .B(_18478_),
    .CI(_18153_),
    .CO(_18479_),
    .S(_18480_));
 FA_X1 _40540_ (.A(_15964_),
    .B(_18481_),
    .CI(_18482_),
    .CO(_16745_),
    .S(_18483_));
 FA_X1 _40541_ (.A(net220),
    .B(net243),
    .CI(_18484_),
    .CO(_18485_),
    .S(_18486_));
 FA_X1 _40542_ (.A(_18487_),
    .B(_18488_),
    .CI(_18489_),
    .CO(_18490_),
    .S(_18491_));
 FA_X1 _40543_ (.A(_18492_),
    .B(_18493_),
    .CI(_18494_),
    .CO(_17992_),
    .S(_18495_));
 FA_X1 _40544_ (.A(_17999_),
    .B(_17245_),
    .CI(_18496_),
    .CO(_18497_),
    .S(_18498_));
 FA_X1 _40545_ (.A(_18499_),
    .B(_18500_),
    .CI(_18501_),
    .CO(_17230_),
    .S(_18502_));
 FA_X1 _40546_ (.A(_18503_),
    .B(_17236_),
    .CI(_18504_),
    .CO(_18505_),
    .S(_18506_));
 FA_X1 _40547_ (.A(_18507_),
    .B(_18508_),
    .CI(_18509_),
    .CO(_18022_),
    .S(_18510_));
 FA_X1 _40548_ (.A(_17212_),
    .B(_18027_),
    .CI(_17217_),
    .CO(_18511_),
    .S(_18512_));
 FA_X1 _40549_ (.A(_18513_),
    .B(_18514_),
    .CI(_18515_),
    .CO(_17172_),
    .S(_18516_));
 FA_X1 _40550_ (.A(_18001_),
    .B(_18006_),
    .CI(_17182_),
    .CO(_18517_),
    .S(_18518_));
 FA_X1 _40551_ (.A(_17153_),
    .B(_18519_),
    .CI(_17144_),
    .CO(_18520_),
    .S(_18521_));
 FA_X1 _40552_ (.A(_17131_),
    .B(_18522_),
    .CI(_18523_),
    .CO(_17620_),
    .S(_18524_));
 FA_X1 _40553_ (.A(_18525_),
    .B(_18526_),
    .CI(_17626_),
    .CO(_18527_),
    .S(_18528_));
 FA_X1 _40554_ (.A(_15651_),
    .B(_18529_),
    .CI(_18530_),
    .CO(_18531_),
    .S(_18532_));
 FA_X1 _40555_ (.A(net172),
    .B(net255),
    .CI(_18533_),
    .CO(_18534_),
    .S(_18535_));
 FA_X1 _40556_ (.A(_18536_),
    .B(_18537_),
    .CI(_18538_),
    .CO(_18539_),
    .S(_18540_));
 FA_X1 _40557_ (.A(_18541_),
    .B(_18542_),
    .CI(_18543_),
    .CO(_18039_),
    .S(_18544_));
 FA_X1 _40558_ (.A(_17107_),
    .B(_18046_),
    .CI(_18545_),
    .CO(_18546_),
    .S(_18547_));
 FA_X1 _40559_ (.A(_18548_),
    .B(_18549_),
    .CI(_18550_),
    .CO(_17092_),
    .S(_18551_));
 FA_X1 _40560_ (.A(_18552_),
    .B(_17098_),
    .CI(_18553_),
    .CO(_18554_),
    .S(_18555_));
 FA_X1 _40561_ (.A(_18556_),
    .B(_18557_),
    .CI(_18558_),
    .CO(_17599_),
    .S(_18559_));
 FA_X1 _40562_ (.A(_18560_),
    .B(_17604_),
    .CI(_17075_),
    .CO(_18561_),
    .S(_18562_));
 FA_X1 _40563_ (.A(_17045_),
    .B(_17583_),
    .CI(_17578_),
    .CO(_18563_),
    .S(_18564_));
 FA_X1 _40564_ (.A(_18565_),
    .B(_18566_),
    .CI(_18567_),
    .CO(_17018_),
    .S(_18568_));
 FA_X1 _40565_ (.A(_17027_),
    .B(_18569_),
    .CI(_18570_),
    .CO(_18067_),
    .S(_18571_));
 FA_X1 _40566_ (.A(_17036_),
    .B(_18572_),
    .CI(_17003_),
    .CO(_18573_),
    .S(_18574_));
 FA_X1 _40567_ (.A(_14944_),
    .B(_18575_),
    .CI(_18576_),
    .CO(_16984_),
    .S(_18577_));
 FA_X1 _40568_ (.A(_18050_),
    .B(_18578_),
    .CI(_18579_),
    .CO(_18580_),
    .S(_18581_));
 FA_X1 _40569_ (.A(net187),
    .B(net267),
    .CI(_18582_),
    .CO(_18583_),
    .S(_18584_));
 FA_X1 _40570_ (.A(_18585_),
    .B(_18586_),
    .CI(_18587_),
    .CO(_18588_),
    .S(_18589_));
 FA_X1 _40571_ (.A(_18240_),
    .B(_16683_),
    .CI(_18590_),
    .CO(_18591_),
    .S(_18592_));
 FA_X1 _40572_ (.A(_18593_),
    .B(_18594_),
    .CI(_18595_),
    .CO(_18229_),
    .S(_18596_));
 FA_X1 _40573_ (.A(_16674_),
    .B(_18597_),
    .CI(_18598_),
    .CO(_18599_),
    .S(_18600_));
 FA_X1 _40574_ (.A(_18601_),
    .B(_18602_),
    .CI(_18603_),
    .CO(_16649_),
    .S(_18604_));
 FA_X1 _40575_ (.A(_16669_),
    .B(_18605_),
    .CI(_17952_),
    .CO(_18606_),
    .S(_18607_));
 FA_X1 _40576_ (.A(_18608_),
    .B(_17938_),
    .CI(_18609_),
    .CO(_17943_),
    .S(_18610_));
 FA_X1 _40577_ (.A(_16617_),
    .B(_17928_),
    .CI(_17948_),
    .CO(_18611_),
    .S(_18612_));
 FA_X1 _40578_ (.A(_18613_),
    .B(_18614_),
    .CI(_18615_),
    .CO(_16594_),
    .S(_18616_));
 FA_X1 _40579_ (.A(net262),
    .B(_16608_),
    .CI(_16599_),
    .CO(_18617_),
    .S(_18618_));
 FA_X1 _40580_ (.A(_18619_),
    .B(_16575_),
    .CI(_16612_),
    .CO(_18620_),
    .S(_18621_));
 FA_X1 _40581_ (.A(_16603_),
    .B(_18622_),
    .CI(_18623_),
    .CO(_18624_),
    .S(_18625_));
 FA_X1 _40582_ (.A(_18626_),
    .B(_18627_),
    .CI(_18624_),
    .CO(_18628_),
    .S(_18629_));
 FA_X1 _40583_ (.A(_18630_),
    .B(_18631_),
    .CI(_18632_),
    .CO(_17650_),
    .S(_18633_));
 FA_X1 _40584_ (.A(net274),
    .B(_18634_),
    .CI(_17642_),
    .CO(_18635_),
    .S(_18636_));
 FA_X1 _40585_ (.A(net211),
    .B(_18637_),
    .CI(_18638_),
    .CO(_18639_),
    .S(_18640_));
 FA_X1 _40586_ (.A(_18641_),
    .B(_18642_),
    .CI(_18643_),
    .CO(_18644_),
    .S(_18645_));
 FA_X1 _40587_ (.A(_18646_),
    .B(_17383_),
    .CI(_17633_),
    .CO(_18647_),
    .S(_18648_));
 FA_X1 _40588_ (.A(_18649_),
    .B(_18650_),
    .CI(_18651_),
    .CO(_17370_),
    .S(_18652_));
 FA_X1 _40589_ (.A(_17292_),
    .B(_18653_),
    .CI(_18654_),
    .CO(_18655_),
    .S(_18656_));
 FA_X1 _40590_ (.A(_18657_),
    .B(_18658_),
    .CI(_18659_),
    .CO(_17267_),
    .S(_18660_));
 FA_X1 _40591_ (.A(_17347_),
    .B(_18661_),
    .CI(_17287_),
    .CO(_18662_),
    .S(_18663_));
 FA_X1 _40592_ (.A(_18664_),
    .B(_18665_),
    .CI(_17310_),
    .CO(_17321_),
    .S(_18666_));
 FA_X1 _40593_ (.A(_17305_),
    .B(_17980_),
    .CI(_17343_),
    .CO(_18667_),
    .S(_18668_));
 FA_X1 _40594_ (.A(_18669_),
    .B(_18670_),
    .CI(_18671_),
    .CO(_17971_),
    .S(_18672_));
 FA_X1 _40595_ (.A(_17420_),
    .B(_18673_),
    .CI(_18674_),
    .CO(_17404_),
    .S(_18675_));
 FA_X1 _40596_ (.A(_18676_),
    .B(_17956_),
    .CI(_17976_),
    .CO(_18677_),
    .S(_18678_));
 FA_X1 _40597_ (.A(_15964_),
    .B(_18679_),
    .CI(_18680_),
    .CO(_17357_),
    .S(_18681_));
 FA_X1 _40598_ (.A(_18682_),
    .B(_18683_),
    .CI(_17387_),
    .CO(_18684_),
    .S(_18685_));
 FA_X1 _40599_ (.A(net149),
    .B(net243),
    .CI(_18686_),
    .CO(_18687_),
    .S(_18688_));
 FA_X1 _40600_ (.A(_18607_),
    .B(_18610_),
    .CI(_16650_),
    .CO(_18689_),
    .S(_18690_));
 FA_X1 _40601_ (.A(_17946_),
    .B(_18606_),
    .CI(_17949_),
    .CO(_18691_),
    .S(_18692_));
 FA_X1 _40602_ (.A(_17945_),
    .B(_18612_),
    .CI(_18616_),
    .CO(_18693_),
    .S(_18694_));
 FA_X1 _40603_ (.A(_16596_),
    .B(_16613_),
    .CI(_18611_),
    .CO(_18695_),
    .S(_18696_));
 FA_X1 _40604_ (.A(_16595_),
    .B(_18621_),
    .CI(_18625_),
    .CO(_18697_),
    .S(_18698_));
 FA_X1 _40605_ (.A(_18633_),
    .B(_18629_),
    .CI(_18620_),
    .CO(_18699_),
    .S(_18700_));
 FA_X1 _40606_ (.A(_17656_),
    .B(_17652_),
    .CI(_18628_),
    .CO(_18701_),
    .S(_18702_));
 FA_X1 _40607_ (.A(_18703_),
    .B(_18704_),
    .CI(_17651_),
    .CO(_18705_),
    .S(_18706_));
 FA_X1 _40608_ (.A(_18707_),
    .B(_18708_),
    .CI(_18709_),
    .CO(_18710_),
    .S(_18711_));
 FA_X1 _40609_ (.A(_18712_),
    .B(_18713_),
    .CI(_18714_),
    .CO(_18715_),
    .S(_18716_));
 FA_X1 _40610_ (.A(_18717_),
    .B(_18718_),
    .CI(_18719_),
    .CO(\g_row[0].g_col[0].mult.stage1.dadda.t1[4] ),
    .S(\g_row[0].g_col[0].mult.stage1.dadda.t2[3] ));
 FA_X1 _40611_ (.A(_18720_),
    .B(_18589_),
    .CI(_18721_),
    .CO(\g_row[0].g_col[0].mult.stage1.dadda.t1[5] ),
    .S(\g_row[0].g_col[0].mult.stage1.dadda.t2[4] ));
 FA_X1 _40612_ (.A(_18722_),
    .B(_16689_),
    .CI(_18723_),
    .CO(_18724_),
    .S(_18725_));
 FA_X1 _40613_ (.A(_18726_),
    .B(_18596_),
    .CI(_16688_),
    .CO(_18727_),
    .S(_18728_));
 FA_X1 _40614_ (.A(_18729_),
    .B(_18231_),
    .CI(_18730_),
    .CO(_18731_),
    .S(_18732_));
 FA_X1 _40615_ (.A(_18230_),
    .B(_18604_),
    .CI(_18600_),
    .CO(_18733_),
    .S(_18734_));
 FA_X1 _40616_ (.A(_18599_),
    .B(_16651_),
    .CI(_16670_),
    .CO(_18735_),
    .S(_18736_));
 FA_X1 _40617_ (.A(_18663_),
    .B(_18666_),
    .CI(_17268_),
    .CO(_18737_),
    .S(_18738_));
 FA_X1 _40618_ (.A(_17323_),
    .B(_17344_),
    .CI(_18662_),
    .CO(_18739_),
    .S(_18740_));
 FA_X1 _40619_ (.A(_17322_),
    .B(_18668_),
    .CI(_18672_),
    .CO(_18741_),
    .S(_18742_));
 FA_X1 _40620_ (.A(_17977_),
    .B(_17973_),
    .CI(_18667_),
    .CO(_18743_),
    .S(_18744_));
 FA_X1 _40621_ (.A(_18678_),
    .B(_18675_),
    .CI(_17972_),
    .CO(_18745_),
    .S(_18746_));
 FA_X1 _40622_ (.A(_17388_),
    .B(_17406_),
    .CI(_18677_),
    .CO(_18747_),
    .S(_18748_));
 FA_X1 _40623_ (.A(_18681_),
    .B(_17405_),
    .CI(_18685_),
    .CO(_18749_),
    .S(_18750_));
 FA_X1 _40624_ (.A(_18751_),
    .B(_18752_),
    .CI(_18684_),
    .CO(_18753_),
    .S(_18754_));
 FA_X1 _40625_ (.A(_18755_),
    .B(_18688_),
    .CI(_17355_),
    .CO(\g_row[0].g_col[1].mult.stage1.dadda.t1[19] ),
    .S(\g_row[0].g_col[1].mult.stage1.dadda.t2[18] ));
 FA_X1 _40626_ (.A(_18756_),
    .B(_18757_),
    .CI(_18758_),
    .CO(_18759_),
    .S(_18760_));
 FA_X1 _40627_ (.A(_18761_),
    .B(_18762_),
    .CI(_18763_),
    .CO(\g_row[0].g_col[1].mult.stage1.dadda.t1[4] ),
    .S(\g_row[0].g_col[1].mult.stage1.dadda.t2[3] ));
 FA_X1 _40628_ (.A(_18764_),
    .B(_18645_),
    .CI(_18765_),
    .CO(\g_row[0].g_col[1].mult.stage1.dadda.t1[5] ),
    .S(\g_row[0].g_col[1].mult.stage1.dadda.t2[4] ));
 FA_X1 _40629_ (.A(_18766_),
    .B(_17639_),
    .CI(_18767_),
    .CO(_18768_),
    .S(_18769_));
 FA_X1 _40630_ (.A(_18770_),
    .B(_18652_),
    .CI(_17638_),
    .CO(_18771_),
    .S(_18772_));
 FA_X1 _40631_ (.A(_17374_),
    .B(_18773_),
    .CI(_18774_),
    .CO(_18775_),
    .S(_18776_));
 FA_X1 _40632_ (.A(_17373_),
    .B(_18660_),
    .CI(_18656_),
    .CO(_18777_),
    .S(_18778_));
 FA_X1 _40633_ (.A(_17269_),
    .B(_17288_),
    .CI(_18655_),
    .CO(_18779_),
    .S(_18780_));
 FA_X1 _40634_ (.A(_18512_),
    .B(_18510_),
    .CI(_17231_),
    .CO(_18781_),
    .S(_18782_));
 FA_X1 _40635_ (.A(_18002_),
    .B(_18024_),
    .CI(_18511_),
    .CO(_18783_),
    .S(_18784_));
 FA_X1 _40636_ (.A(_18516_),
    .B(_18518_),
    .CI(_18023_),
    .CO(_18785_),
    .S(_18786_));
 FA_X1 _40637_ (.A(_17145_),
    .B(_17174_),
    .CI(_18517_),
    .CO(_18787_),
    .S(_18788_));
 FA_X1 _40638_ (.A(_17173_),
    .B(_18524_),
    .CI(_18521_),
    .CO(_18789_),
    .S(_18790_));
 FA_X1 _40639_ (.A(_17627_),
    .B(_17622_),
    .CI(_18520_),
    .CO(_18791_),
    .S(_18792_));
 FA_X1 _40640_ (.A(_18528_),
    .B(_18532_),
    .CI(_17621_),
    .CO(_18793_),
    .S(_18794_));
 FA_X1 _40641_ (.A(_18795_),
    .B(_18796_),
    .CI(_18527_),
    .CO(_18797_),
    .S(_18798_));
 FA_X1 _40642_ (.A(_18799_),
    .B(_18800_),
    .CI(_18801_),
    .CO(_18802_),
    .S(_18803_));
 FA_X1 _40643_ (.A(_18804_),
    .B(_18805_),
    .CI(_18806_),
    .CO(_18807_),
    .S(_18808_));
 FA_X1 _40644_ (.A(_18809_),
    .B(_18810_),
    .CI(_18811_),
    .CO(\g_row[0].g_col[2].mult.stage1.dadda.t1[4] ),
    .S(\g_row[0].g_col[2].mult.stage1.dadda.t2[3] ));
 FA_X1 _40645_ (.A(_18812_),
    .B(_18491_),
    .CI(_18813_),
    .CO(\g_row[0].g_col[2].mult.stage1.dadda.t1[5] ),
    .S(\g_row[0].g_col[2].mult.stage1.dadda.t2[4] ));
 FA_X1 _40646_ (.A(_18814_),
    .B(_17251_),
    .CI(_18815_),
    .CO(_18816_),
    .S(_18817_));
 FA_X1 _40647_ (.A(_18819_),
    .B(_18495_),
    .CI(_17250_),
    .CO(_18820_),
    .S(_18821_));
 FA_X1 _40648_ (.A(_18822_),
    .B(_17994_),
    .CI(_18823_),
    .CO(_18824_),
    .S(_18825_));
 FA_X1 _40649_ (.A(_18502_),
    .B(_18506_),
    .CI(_17993_),
    .CO(_18826_),
    .S(_18827_));
 FA_X1 _40650_ (.A(_17213_),
    .B(_17232_),
    .CI(_18505_),
    .CO(_18828_),
    .S(_18829_));
 FA_X1 _40651_ (.A(_17093_),
    .B(_18559_),
    .CI(_18562_),
    .CO(_18830_),
    .S(_18831_));
 FA_X1 _40652_ (.A(_17579_),
    .B(_17601_),
    .CI(_18561_),
    .CO(_18832_),
    .S(_18833_));
 FA_X1 _40653_ (.A(_18568_),
    .B(_18564_),
    .CI(_17600_),
    .CO(_18834_),
    .S(_18835_));
 FA_X1 _40654_ (.A(_17020_),
    .B(_17037_),
    .CI(_18563_),
    .CO(_18836_),
    .S(_18837_));
 FA_X1 _40655_ (.A(_17019_),
    .B(_18571_),
    .CI(_18574_),
    .CO(_18838_),
    .S(_18839_));
 FA_X1 _40656_ (.A(_18051_),
    .B(_18069_),
    .CI(_18573_),
    .CO(_18840_),
    .S(_18841_));
 FA_X1 _40657_ (.A(_18581_),
    .B(_18577_),
    .CI(_18068_),
    .CO(_18842_),
    .S(_18843_));
 FA_X1 _40658_ (.A(_18844_),
    .B(_18845_),
    .CI(_18580_),
    .CO(_18846_),
    .S(_18847_));
 FA_X1 _40659_ (.A(_16982_),
    .B(_18584_),
    .CI(_18848_),
    .CO(\g_row[0].g_col[3].mult.stage1.dadda.t1[19] ),
    .S(\g_row[0].g_col[3].mult.stage1.dadda.t2[18] ));
 FA_X1 _40660_ (.A(_18849_),
    .B(_18850_),
    .CI(_18851_),
    .CO(_18852_),
    .S(_18853_));
 FA_X1 _40661_ (.A(_18854_),
    .B(_18855_),
    .CI(_18856_),
    .CO(\g_row[0].g_col[3].mult.stage1.dadda.t1[4] ),
    .S(\g_row[0].g_col[3].mult.stage1.dadda.t2[3] ));
 FA_X1 _40662_ (.A(_18857_),
    .B(_18540_),
    .CI(_18858_),
    .CO(\g_row[0].g_col[3].mult.stage1.dadda.t1[5] ),
    .S(\g_row[0].g_col[3].mult.stage1.dadda.t2[4] ));
 FA_X1 _40663_ (.A(_18859_),
    .B(_18860_),
    .CI(_17113_),
    .CO(_18861_),
    .S(_18862_));
 FA_X1 _40664_ (.A(_17112_),
    .B(_18544_),
    .CI(_18864_),
    .CO(_18865_),
    .S(_18866_));
 FA_X1 _40665_ (.A(_18867_),
    .B(_18041_),
    .CI(_18868_),
    .CO(_18869_),
    .S(_18870_));
 FA_X1 _40666_ (.A(_18551_),
    .B(_18555_),
    .CI(_18040_),
    .CO(_18871_),
    .S(_18872_));
 FA_X1 _40667_ (.A(_17076_),
    .B(_17094_),
    .CI(_18554_),
    .CO(_18873_),
    .S(_18874_));
 FA_X1 _40668_ (.A(_16921_),
    .B(_16943_),
    .CI(_18385_),
    .CO(_18875_),
    .S(_18876_));
 FA_X1 _40669_ (.A(_18396_),
    .B(_18399_),
    .CI(_16920_),
    .CO(_18877_),
    .S(_18878_));
 FA_X1 _40670_ (.A(_18405_),
    .B(_18401_),
    .CI(_18395_),
    .CO(_18879_),
    .S(_18880_));
 FA_X1 _40671_ (.A(_18101_),
    .B(_18105_),
    .CI(_18400_),
    .CO(_18881_),
    .S(_18882_));
 FA_X1 _40672_ (.A(_18408_),
    .B(_18411_),
    .CI(_18100_),
    .CO(_18883_),
    .S(_18884_));
 FA_X1 _40673_ (.A(_16870_),
    .B(_16879_),
    .CI(_18410_),
    .CO(_18885_),
    .S(_18886_));
 FA_X1 _40674_ (.A(_16869_),
    .B(_18419_),
    .CI(_18415_),
    .CO(_18887_),
    .S(_18888_));
 FA_X1 _40675_ (.A(_18889_),
    .B(_18414_),
    .CI(_18890_),
    .CO(_18891_),
    .S(_18892_));
 FA_X1 _40676_ (.A(_18893_),
    .B(_18894_),
    .CI(_18895_),
    .CO(_18896_),
    .S(_18897_));
 FA_X1 _40677_ (.A(_18898_),
    .B(_18713_),
    .CI(_18899_),
    .CO(_18900_),
    .S(_18901_));
 FA_X1 _40678_ (.A(_18902_),
    .B(_18903_),
    .CI(_18904_),
    .CO(\g_row[1].g_col[0].mult.stage1.dadda.t1[4] ),
    .S(\g_row[1].g_col[0].mult.stage1.dadda.t2[3] ));
 FA_X1 _40679_ (.A(_18905_),
    .B(_18906_),
    .CI(_18076_),
    .CO(\g_row[1].g_col[0].mult.stage1.dadda.t1[5] ),
    .S(\g_row[1].g_col[0].mult.stage1.dadda.t2[4] ));
 FA_X1 _40680_ (.A(_18907_),
    .B(_18908_),
    .CI(_18375_),
    .CO(_18909_),
    .S(_18910_));
 FA_X1 _40681_ (.A(_16970_),
    .B(_18911_),
    .CI(_18374_),
    .CO(_18912_),
    .S(_18913_));
 FA_X1 _40682_ (.A(_18379_),
    .B(_18914_),
    .CI(_18915_),
    .CO(_18916_),
    .S(_18917_));
 FA_X1 _40683_ (.A(_17570_),
    .B(_17565_),
    .CI(_18378_),
    .CO(_18918_),
    .S(_18919_));
 FA_X1 _40684_ (.A(_18386_),
    .B(_17564_),
    .CI(_18389_),
    .CO(_18920_),
    .S(_18921_));
 FA_X1 _40685_ (.A(_18461_),
    .B(_18464_),
    .CI(_18453_),
    .CO(_18922_),
    .S(_18923_));
 FA_X1 _40686_ (.A(_17533_),
    .B(_17529_),
    .CI(_18460_),
    .CO(_18924_),
    .S(_18925_));
 FA_X1 _40687_ (.A(_18470_),
    .B(_18466_),
    .CI(_17528_),
    .CO(_18926_),
    .S(_18927_));
 FA_X1 _40688_ (.A(_16781_),
    .B(_16798_),
    .CI(_18465_),
    .CO(_18928_),
    .S(_18929_));
 FA_X1 _40689_ (.A(_18473_),
    .B(_18476_),
    .CI(_16780_),
    .CO(_18930_),
    .S(_18931_));
 FA_X1 _40690_ (.A(_18149_),
    .B(_18154_),
    .CI(_18472_),
    .CO(_18932_),
    .S(_18933_));
 FA_X1 _40691_ (.A(_18148_),
    .B(_18483_),
    .CI(_18480_),
    .CO(_18934_),
    .S(_18935_));
 FA_X1 _40692_ (.A(_18936_),
    .B(_18937_),
    .CI(_18479_),
    .CO(_18938_),
    .S(_18939_));
 FA_X1 _40693_ (.A(_18940_),
    .B(_18941_),
    .CI(_18942_),
    .CO(_18943_),
    .S(_18944_));
 FA_X1 _40694_ (.A(_18945_),
    .B(_18757_),
    .CI(_18946_),
    .CO(_18947_),
    .S(_18948_));
 FA_X1 _40695_ (.A(_18949_),
    .B(_18950_),
    .CI(_18951_),
    .CO(\g_row[1].g_col[1].mult.stage1.dadda.t1[4] ),
    .S(\g_row[1].g_col[1].mult.stage1.dadda.t2[3] ));
 FA_X1 _40696_ (.A(_18952_),
    .B(_18953_),
    .CI(_18427_),
    .CO(\g_row[1].g_col[1].mult.stage1.dadda.t1[5] ),
    .S(\g_row[1].g_col[1].mult.stage1.dadda.t2[4] ));
 FA_X1 _40697_ (.A(_18131_),
    .B(_18954_),
    .CI(_18955_),
    .CO(_18956_),
    .S(_18957_));
 FA_X1 _40698_ (.A(_18130_),
    .B(_18958_),
    .CI(_18440_),
    .CO(_18959_),
    .S(_18960_));
 FA_X1 _40699_ (.A(_18448_),
    .B(_18444_),
    .CI(_18961_),
    .CO(_18962_),
    .S(_18963_));
 FA_X1 _40700_ (.A(_16832_),
    .B(_16847_),
    .CI(_18443_),
    .CO(_18964_),
    .S(_18965_));
 FA_X1 _40701_ (.A(_18458_),
    .B(_18454_),
    .CI(_16831_),
    .CO(_18966_),
    .S(_18967_));
 FA_X1 _40702_ (.A(_17887_),
    .B(_17883_),
    .CI(_18291_),
    .CO(_18968_),
    .S(_18969_));
 FA_X1 _40703_ (.A(_17882_),
    .B(_18300_),
    .CI(_18297_),
    .CO(_18970_),
    .S(_18971_));
 FA_X1 _40704_ (.A(_17469_),
    .B(_17490_),
    .CI(_18296_),
    .CO(_18972_),
    .S(_18973_));
 FA_X1 _40705_ (.A(_18302_),
    .B(_18305_),
    .CI(_17468_),
    .CO(_18974_),
    .S(_18975_));
 FA_X1 _40706_ (.A(_17837_),
    .B(_17856_),
    .CI(_18301_),
    .CO(_18976_),
    .S(_18977_));
 FA_X1 _40707_ (.A(_17855_),
    .B(_18309_),
    .CI(_18313_),
    .CO(_18978_),
    .S(_18979_));
 FA_X1 _40708_ (.A(_18178_),
    .B(_18191_),
    .CI(_18312_),
    .CO(_18980_),
    .S(_18981_));
 FA_X1 _40709_ (.A(_18982_),
    .B(_18983_),
    .CI(_18190_),
    .CO(_18984_),
    .S(_18985_));
 FA_X1 _40710_ (.A(_18986_),
    .B(_17823_),
    .CI(_18320_),
    .CO(\g_row[1].g_col[2].mult.stage1.dadda.t1[19] ),
    .S(\g_row[1].g_col[2].mult.stage1.dadda.t2[18] ));
 FA_X1 _40711_ (.A(_18987_),
    .B(_18805_),
    .CI(_18988_),
    .CO(_18989_),
    .S(_18990_));
 FA_X1 _40712_ (.A(_18991_),
    .B(_18992_),
    .CI(_18993_),
    .CO(\g_row[1].g_col[2].mult.stage1.dadda.t1[4] ),
    .S(\g_row[1].g_col[2].mult.stage1.dadda.t2[3] ));
 FA_X1 _40713_ (.A(_17430_),
    .B(_18994_),
    .CI(_18995_),
    .CO(\g_row[1].g_col[2].mult.stage1.dadda.t1[5] ),
    .S(\g_row[1].g_col[2].mult.stage1.dadda.t2[4] ));
 FA_X1 _40714_ (.A(_18281_),
    .B(_18996_),
    .CI(_18997_),
    .CO(_18998_),
    .S(_18999_));
 FA_X1 _40715_ (.A(_18280_),
    .B(_19000_),
    .CI(_18170_),
    .CO(_19001_),
    .S(_19002_));
 FA_X1 _40716_ (.A(_18289_),
    .B(_18285_),
    .CI(_19003_),
    .CO(_19004_),
    .S(_19005_));
 FA_X1 _40717_ (.A(_18284_),
    .B(_17914_),
    .CI(_17919_),
    .CO(_19006_),
    .S(_19007_));
 FA_X1 _40718_ (.A(_18292_),
    .B(_18295_),
    .CI(_17913_),
    .CO(_19008_),
    .S(_19009_));
 FA_X1 _40719_ (.A(_18348_),
    .B(_18345_),
    .CI(_18216_),
    .CO(_19010_),
    .S(_19011_));
 FA_X1 _40720_ (.A(_17756_),
    .B(_17778_),
    .CI(_18347_),
    .CO(_19012_),
    .S(_19013_));
 FA_X1 _40721_ (.A(_18352_),
    .B(_17777_),
    .CI(_18354_),
    .CO(_19014_),
    .S(_19015_));
 FA_X1 _40722_ (.A(_17732_),
    .B(_17703_),
    .CI(_18353_),
    .CO(_19016_),
    .S(_19017_));
 FA_X1 _40723_ (.A(_18360_),
    .B(_18357_),
    .CI(_17731_),
    .CO(_19018_),
    .S(_19019_));
 FA_X1 _40724_ (.A(_18274_),
    .B(_18256_),
    .CI(_18359_),
    .CO(_19020_),
    .S(_19021_));
 FA_X1 _40725_ (.A(_18363_),
    .B(_18367_),
    .CI(_18273_),
    .CO(_19022_),
    .S(_19023_));
 FA_X1 _40726_ (.A(_18366_),
    .B(_19024_),
    .CI(_19025_),
    .CO(_19026_),
    .S(_19027_));
 FA_X1 _40727_ (.A(_18370_),
    .B(_19028_),
    .CI(_17677_),
    .CO(\g_row[1].g_col[3].mult.stage1.dadda.t1[19] ),
    .S(\g_row[1].g_col[3].mult.stage1.dadda.t2[18] ));
 FA_X1 _40728_ (.A(_19029_),
    .B(_18850_),
    .CI(_19030_),
    .CO(_19031_),
    .S(_19032_));
 FA_X1 _40729_ (.A(_19033_),
    .B(_19034_),
    .CI(_19035_),
    .CO(\g_row[1].g_col[3].mult.stage1.dadda.t1[4] ),
    .S(\g_row[1].g_col[3].mult.stage1.dadda.t2[3] ));
 FA_X1 _40730_ (.A(_19036_),
    .B(_19037_),
    .CI(_18326_),
    .CO(\g_row[1].g_col[3].mult.stage1.dadda.t1[5] ),
    .S(\g_row[1].g_col[3].mult.stage1.dadda.t2[4] ));
 FA_X1 _40731_ (.A(_17440_),
    .B(_19038_),
    .CI(_19039_),
    .CO(_19040_),
    .S(_19041_));
 FA_X1 _40732_ (.A(_18330_),
    .B(_19042_),
    .CI(_17439_),
    .CO(_19043_),
    .S(_19044_));
 FA_X1 _40733_ (.A(_19045_),
    .B(_19046_),
    .CI(_17815_),
    .CO(_19047_),
    .S(_19048_));
 FA_X1 _40734_ (.A(_17814_),
    .B(_18337_),
    .CI(_18341_),
    .CO(_19049_),
    .S(_19050_));
 FA_X1 _40735_ (.A(_18199_),
    .B(_18217_),
    .CI(_18340_),
    .CO(_19051_),
    .S(_19052_));
 FA_X1 _40736_ (.A(_14989_),
    .B(_14995_),
    .CI(_14558_),
    .CO(_19053_),
    .S(_19054_));
 FA_X1 _40737_ (.A(_14994_),
    .B(_15345_),
    .CI(_15343_),
    .CO(_19055_),
    .S(_19056_));
 FA_X1 _40738_ (.A(_15337_),
    .B(_15333_),
    .CI(_15344_),
    .CO(_19057_),
    .S(_19058_));
 FA_X1 _40739_ (.A(_15299_),
    .B(_15295_),
    .CI(_15336_),
    .CO(_19059_),
    .S(_19060_));
 FA_X1 _40740_ (.A(_15272_),
    .B(_15267_),
    .CI(_15298_),
    .CO(_19061_),
    .S(_19062_));
 FA_X1 _40741_ (.A(_15226_),
    .B(_15221_),
    .CI(_15271_),
    .CO(_19063_),
    .S(_19064_));
 FA_X1 _40742_ (.A(_15204_),
    .B(_15199_),
    .CI(_15225_),
    .CO(_19065_),
    .S(_19066_));
 FA_X1 _40743_ (.A(_19067_),
    .B(_19068_),
    .CI(_15203_),
    .CO(_19069_),
    .S(_19070_));
 FA_X1 _40744_ (.A(_15162_),
    .B(_19071_),
    .CI(_15127_),
    .CO(\g_row[2].g_col[0].mult.stage1.dadda.t1[19] ),
    .S(\g_row[2].g_col[0].mult.stage1.dadda.t2[18] ));
 FA_X1 _40745_ (.A(_19072_),
    .B(_18713_),
    .CI(_19073_),
    .CO(_19074_),
    .S(_19075_));
 FA_X1 _40746_ (.A(_19076_),
    .B(_19077_),
    .CI(_19078_),
    .CO(_19079_),
    .S(_19080_));
 FA_X1 _40747_ (.A(_19081_),
    .B(_14637_),
    .CI(_19082_),
    .CO(\g_row[2].g_col[0].mult.stage1.dadda.t1[5] ),
    .S(\g_row[2].g_col[0].mult.stage1.dadda.t2[4] ));
 FA_X1 _40748_ (.A(_19083_),
    .B(_14632_),
    .CI(_19084_),
    .CO(_19085_),
    .S(_19086_));
 FA_X1 _40749_ (.A(_14619_),
    .B(_19088_),
    .CI(_14631_),
    .CO(_19089_),
    .S(_19090_));
 FA_X1 _40750_ (.A(_19091_),
    .B(_14607_),
    .CI(_19092_),
    .CO(_19093_),
    .S(_19094_));
 FA_X1 _40751_ (.A(_14593_),
    .B(_14589_),
    .CI(_14606_),
    .CO(_19095_),
    .S(_19096_));
 FA_X1 _40752_ (.A(_14592_),
    .B(_14540_),
    .CI(_14559_),
    .CO(_19097_),
    .S(_19098_));
 FA_X1 _40753_ (.A(_16141_),
    .B(_16144_),
    .CI(_16161_),
    .CO(_19099_),
    .S(_19100_));
 FA_X1 _40754_ (.A(_16119_),
    .B(_16116_),
    .CI(_16140_),
    .CO(_19101_),
    .S(_19102_));
 FA_X1 _40755_ (.A(_16095_),
    .B(_16091_),
    .CI(_16115_),
    .CO(_19103_),
    .S(_19104_));
 FA_X1 _40756_ (.A(_16067_),
    .B(_16064_),
    .CI(_16090_),
    .CO(_19105_),
    .S(_19106_));
 FA_X1 _40757_ (.A(_16040_),
    .B(_16037_),
    .CI(_16063_),
    .CO(_19107_),
    .S(_19108_));
 FA_X1 _40758_ (.A(_16004_),
    .B(_16013_),
    .CI(_16036_),
    .CO(_19109_),
    .S(_19110_));
 FA_X1 _40759_ (.A(_16513_),
    .B(_16517_),
    .CI(_16003_),
    .CO(_19111_),
    .S(_19112_));
 FA_X1 _40760_ (.A(_19113_),
    .B(_19114_),
    .CI(_16512_),
    .CO(_19115_),
    .S(_19116_));
 FA_X1 _40761_ (.A(_19117_),
    .B(_19118_),
    .CI(_19119_),
    .CO(_19120_),
    .S(_19121_));
 FA_X1 _40762_ (.A(_19122_),
    .B(_18757_),
    .CI(_19123_),
    .CO(_19124_),
    .S(_19125_));
 FA_X1 _40763_ (.A(_19126_),
    .B(_19127_),
    .CI(_19128_),
    .CO(\g_row[2].g_col[1].mult.stage1.dadda.t1[4] ),
    .S(\g_row[2].g_col[1].mult.stage1.dadda.t2[3] ));
 FA_X1 _40764_ (.A(_16223_),
    .B(_19129_),
    .CI(_19130_),
    .CO(\g_row[2].g_col[1].mult.stage1.dadda.t1[5] ),
    .S(\g_row[2].g_col[1].mult.stage1.dadda.t2[4] ));
 FA_X1 _40765_ (.A(_19131_),
    .B(_16218_),
    .CI(_19132_),
    .CO(_19133_),
    .S(_19134_));
 FA_X1 _40766_ (.A(_16209_),
    .B(_19135_),
    .CI(_16217_),
    .CO(_19136_),
    .S(_19137_));
 FA_X1 _40767_ (.A(_19138_),
    .B(_16192_),
    .CI(_19139_),
    .CO(_19140_),
    .S(_19141_));
 FA_X1 _40768_ (.A(_16178_),
    .B(_16182_),
    .CI(_16191_),
    .CO(_19142_),
    .S(_19143_));
 FA_X1 _40769_ (.A(_16177_),
    .B(_16162_),
    .CI(_16165_),
    .CO(_19144_),
    .S(_19145_));
 FA_X1 _40770_ (.A(_16713_),
    .B(_16693_),
    .CI(_16696_),
    .CO(_19146_),
    .S(_19147_));
 FA_X1 _40771_ (.A(_14663_),
    .B(_14685_),
    .CI(_16692_),
    .CO(_19148_),
    .S(_19149_));
 FA_X1 _40772_ (.A(_15133_),
    .B(_15154_),
    .CI(_14662_),
    .CO(_19150_),
    .S(_19151_));
 FA_X1 _40773_ (.A(_15411_),
    .B(_15429_),
    .CI(_15132_),
    .CO(_19152_),
    .S(_19153_));
 FA_X1 _40774_ (.A(_15699_),
    .B(_15704_),
    .CI(_15410_),
    .CO(_19154_),
    .S(_19155_));
 FA_X1 _40775_ (.A(_15762_),
    .B(_15770_),
    .CI(_15703_),
    .CO(_19156_),
    .S(_19157_));
 FA_X1 _40776_ (.A(_16476_),
    .B(_16484_),
    .CI(_15769_),
    .CO(_19158_),
    .S(_19159_));
 FA_X1 _40777_ (.A(_19160_),
    .B(_19161_),
    .CI(_16483_),
    .CO(_19162_),
    .S(_19163_));
 FA_X1 _40778_ (.A(_19164_),
    .B(_15707_),
    .CI(_16728_),
    .CO(\g_row[2].g_col[2].mult.stage1.dadda.t1[19] ),
    .S(\g_row[2].g_col[2].mult.stage1.dadda.t2[18] ));
 FA_X1 _40779_ (.A(_19165_),
    .B(_18805_),
    .CI(_19166_),
    .CO(_19167_),
    .S(_19168_));
 FA_X1 _40780_ (.A(_19169_),
    .B(_19170_),
    .CI(_19171_),
    .CO(_19172_),
    .S(_19173_));
 FA_X1 _40781_ (.A(_16564_),
    .B(_19174_),
    .CI(_19175_),
    .CO(\g_row[2].g_col[2].mult.stage1.dadda.t1[5] ),
    .S(\g_row[2].g_col[2].mult.stage1.dadda.t2[4] ));
 FA_X1 _40782_ (.A(_19176_),
    .B(_16559_),
    .CI(_19177_),
    .CO(_19178_),
    .S(_19179_));
 FA_X1 _40783_ (.A(_19180_),
    .B(_16550_),
    .CI(_16558_),
    .CO(_19181_),
    .S(_19182_));
 FA_X1 _40784_ (.A(_16537_),
    .B(_16527_),
    .CI(_19183_),
    .CO(_19184_),
    .S(_19185_));
 FA_X1 _40785_ (.A(_16526_),
    .B(_16736_),
    .CI(_16732_),
    .CO(_19186_),
    .S(_19187_));
 FA_X1 _40786_ (.A(_16714_),
    .B(_16731_),
    .CI(_16717_),
    .CO(_19188_),
    .S(_19189_));
 FA_X1 _40787_ (.A(_15070_),
    .B(_15048_),
    .CI(_15012_),
    .CO(_19190_),
    .S(_19191_));
 FA_X1 _40788_ (.A(_15076_),
    .B(_15097_),
    .CI(_15047_),
    .CO(_19192_),
    .S(_19193_));
 FA_X1 _40789_ (.A(_15075_),
    .B(_15103_),
    .CI(_15124_),
    .CO(_19194_),
    .S(_19195_));
 FA_X1 _40790_ (.A(_15188_),
    .B(_15195_),
    .CI(_15102_),
    .CO(_19196_),
    .S(_19197_));
 FA_X1 _40791_ (.A(_15259_),
    .B(_15264_),
    .CI(_15194_),
    .CO(_19198_),
    .S(_19199_));
 FA_X1 _40792_ (.A(_15321_),
    .B(_15329_),
    .CI(_15263_),
    .CO(_19200_),
    .S(_19201_));
 FA_X1 _40793_ (.A(_15348_),
    .B(_15352_),
    .CI(_15328_),
    .CO(_19202_),
    .S(_19203_));
 FA_X1 _40794_ (.A(_19204_),
    .B(_19205_),
    .CI(_15351_),
    .CO(_19206_),
    .S(_19207_));
 FA_X1 _40795_ (.A(_19208_),
    .B(_14615_),
    .CI(_14576_),
    .CO(\g_row[2].g_col[3].mult.stage1.dadda.t1[19] ),
    .S(\g_row[2].g_col[3].mult.stage1.dadda.t2[18] ));
 FA_X1 _40796_ (.A(_19209_),
    .B(_18850_),
    .CI(_19210_),
    .CO(_19211_),
    .S(_19212_));
 FA_X1 _40797_ (.A(_19213_),
    .B(_19214_),
    .CI(_19215_),
    .CO(_19216_),
    .S(_19217_));
 FA_X1 _40798_ (.A(_19218_),
    .B(_15372_),
    .CI(_19219_),
    .CO(\g_row[2].g_col[3].mult.stage1.dadda.t1[5] ),
    .S(\g_row[2].g_col[3].mult.stage1.dadda.t2[4] ));
 FA_X1 _40799_ (.A(_15487_),
    .B(_19220_),
    .CI(_19221_),
    .CO(_19222_),
    .S(_19223_));
 FA_X1 _40800_ (.A(_19224_),
    .B(_15607_),
    .CI(_15486_),
    .CO(_19225_),
    .S(_19226_));
 FA_X1 _40801_ (.A(_15671_),
    .B(_15676_),
    .CI(_19227_),
    .CO(_19228_),
    .S(_19229_));
 FA_X1 _40802_ (.A(_15670_),
    .B(_15686_),
    .CI(_15682_),
    .CO(_19230_),
    .S(_19231_));
 FA_X1 _40803_ (.A(_15013_),
    .B(_15032_),
    .CI(_15681_),
    .CO(_19232_),
    .S(_19233_));
 FA_X1 _40804_ (.A(_16341_),
    .B(_16347_),
    .CI(_16318_),
    .CO(_19234_),
    .S(_19235_));
 FA_X1 _40805_ (.A(_16346_),
    .B(_16368_),
    .CI(_16375_),
    .CO(_19236_),
    .S(_19237_));
 FA_X1 _40806_ (.A(_16401_),
    .B(_16396_),
    .CI(_16374_),
    .CO(_19238_),
    .S(_19239_));
 FA_X1 _40807_ (.A(_16408_),
    .B(_16400_),
    .CI(_16425_),
    .CO(_19240_),
    .S(_19241_));
 FA_X1 _40808_ (.A(_16430_),
    .B(_16443_),
    .CI(_16407_),
    .CO(_19242_),
    .S(_19243_));
 FA_X1 _40809_ (.A(_16451_),
    .B(_16460_),
    .CI(_16429_),
    .CO(_19244_),
    .S(_19245_));
 FA_X1 _40810_ (.A(_16464_),
    .B(_16472_),
    .CI(_16450_),
    .CO(_19246_),
    .S(_19247_));
 FA_X1 _40811_ (.A(_19248_),
    .B(_19249_),
    .CI(_16471_),
    .CO(_19250_),
    .S(_19251_));
 FA_X1 _40812_ (.A(_16491_),
    .B(_19252_),
    .CI(_16495_),
    .CO(\g_row[3].g_col[0].mult.stage1.dadda.t1[19] ),
    .S(\g_row[3].g_col[0].mult.stage1.dadda.t2[18] ));
 FA_X1 _40813_ (.A(_19253_),
    .B(_18713_),
    .CI(_19254_),
    .CO(_19255_),
    .S(_19256_));
 FA_X1 _40814_ (.A(_19257_),
    .B(_19258_),
    .CI(_19259_),
    .CO(_19260_),
    .S(_19261_));
 FA_X1 _40815_ (.A(_16228_),
    .B(_19262_),
    .CI(_19263_),
    .CO(\g_row[3].g_col[0].mult.stage1.dadda.t1[5] ),
    .S(\g_row[3].g_col[0].mult.stage1.dadda.t2[4] ));
 FA_X1 _40816_ (.A(_19264_),
    .B(_16238_),
    .CI(_19265_),
    .CO(_19266_),
    .S(_19267_));
 FA_X1 _40817_ (.A(_16237_),
    .B(_16243_),
    .CI(_19269_),
    .CO(_19270_),
    .S(_19271_));
 FA_X1 _40818_ (.A(_19272_),
    .B(_19273_),
    .CI(_16269_),
    .CO(_19274_),
    .S(_19275_));
 FA_X1 _40819_ (.A(_16293_),
    .B(_16284_),
    .CI(_16268_),
    .CO(_19276_),
    .S(_19277_));
 FA_X1 _40820_ (.A(_16312_),
    .B(_16319_),
    .CI(_16292_),
    .CO(_19278_),
    .S(_19279_));
 FA_X1 _40821_ (.A(_15826_),
    .B(_15848_),
    .CI(_15799_),
    .CO(_19280_),
    .S(_19281_));
 FA_X1 _40822_ (.A(_15855_),
    .B(_15877_),
    .CI(_15825_),
    .CO(_19282_),
    .S(_19283_));
 FA_X1 _40823_ (.A(_15882_),
    .B(_15903_),
    .CI(_15854_),
    .CO(_19284_),
    .S(_19285_));
 FA_X1 _40824_ (.A(_15910_),
    .B(_15928_),
    .CI(_15881_),
    .CO(_19286_),
    .S(_19287_));
 FA_X1 _40825_ (.A(_15941_),
    .B(_15946_),
    .CI(_15909_),
    .CO(_19288_),
    .S(_19289_));
 FA_X1 _40826_ (.A(_15963_),
    .B(_15955_),
    .CI(_15945_),
    .CO(_19290_),
    .S(_19291_));
 FA_X1 _40827_ (.A(_15968_),
    .B(_15962_),
    .CI(_15976_),
    .CO(_19292_),
    .S(_19293_));
 FA_X1 _40828_ (.A(_15975_),
    .B(_19294_),
    .CI(_19295_),
    .CO(_19296_),
    .S(_19297_));
 FA_X1 _40829_ (.A(_19298_),
    .B(_19299_),
    .CI(_19300_),
    .CO(_19301_),
    .S(_19302_));
 FA_X1 _40830_ (.A(_19303_),
    .B(_18757_),
    .CI(_19304_),
    .CO(_19305_),
    .S(_19306_));
 FA_X1 _40831_ (.A(_19307_),
    .B(_19308_),
    .CI(_19309_),
    .CO(_19310_),
    .S(_19311_));
 FA_X1 _40832_ (.A(_19312_),
    .B(_15712_),
    .CI(_19313_),
    .CO(\g_row[3].g_col[1].mult.stage1.dadda.t1[5] ),
    .S(\g_row[3].g_col[1].mult.stage1.dadda.t2[4] ));
 FA_X1 _40833_ (.A(_15722_),
    .B(_19314_),
    .CI(_19315_),
    .CO(_19316_),
    .S(_19317_));
 FA_X1 _40834_ (.A(_19319_),
    .B(_15735_),
    .CI(_15721_),
    .CO(_19320_),
    .S(_19321_));
 FA_X1 _40835_ (.A(_15744_),
    .B(_19322_),
    .CI(_19323_),
    .CO(_19324_),
    .S(_19325_));
 FA_X1 _40836_ (.A(_15794_),
    .B(_15779_),
    .CI(_15743_),
    .CO(_19326_),
    .S(_19327_));
 FA_X1 _40837_ (.A(_15800_),
    .B(_15778_),
    .CI(_15819_),
    .CO(_19328_),
    .S(_19329_));
 FA_X1 _40838_ (.A(_15494_),
    .B(_15516_),
    .CI(_15457_),
    .CO(_19330_),
    .S(_19331_));
 FA_X1 _40839_ (.A(_15522_),
    .B(_15543_),
    .CI(_15493_),
    .CO(_19332_),
    .S(_19333_));
 FA_X1 _40840_ (.A(_15549_),
    .B(_15570_),
    .CI(_15521_),
    .CO(_19334_),
    .S(_19335_));
 FA_X1 _40841_ (.A(_15577_),
    .B(_15594_),
    .CI(_15548_),
    .CO(_19336_),
    .S(_19337_));
 FA_X1 _40842_ (.A(_15612_),
    .B(_15576_),
    .CI(_15625_),
    .CO(_19338_),
    .S(_19339_));
 FA_X1 _40843_ (.A(_15633_),
    .B(_15611_),
    .CI(_15642_),
    .CO(_19340_),
    .S(_19341_));
 FA_X1 _40844_ (.A(_15650_),
    .B(_15655_),
    .CI(_15632_),
    .CO(_19342_),
    .S(_19343_));
 FA_X1 _40845_ (.A(_19344_),
    .B(_19345_),
    .CI(_15649_),
    .CO(_19346_),
    .S(_19347_));
 FA_X1 _40846_ (.A(_19348_),
    .B(_19349_),
    .CI(_19350_),
    .CO(_19351_),
    .S(_19352_));
 FA_X1 _40847_ (.A(_19353_),
    .B(_18805_),
    .CI(_19354_),
    .CO(_19355_),
    .S(_19356_));
 FA_X1 _40848_ (.A(_19357_),
    .B(_19358_),
    .CI(_19359_),
    .CO(_19360_),
    .S(_19361_));
 FA_X1 _40849_ (.A(_15357_),
    .B(_19362_),
    .CI(_19363_),
    .CO(\g_row[3].g_col[2].mult.stage1.dadda.t1[5] ),
    .S(\g_row[3].g_col[2].mult.stage1.dadda.t2[4] ));
 FA_X1 _40850_ (.A(_15367_),
    .B(_19364_),
    .CI(_19365_),
    .CO(_19366_),
    .S(_19367_));
 FA_X1 _40851_ (.A(_15385_),
    .B(_19368_),
    .CI(_15366_),
    .CO(_19369_),
    .S(_19370_));
 FA_X1 _40852_ (.A(_19371_),
    .B(_15394_),
    .CI(_15404_),
    .CO(_19372_),
    .S(_19373_));
 FA_X1 _40853_ (.A(_15437_),
    .B(_15452_),
    .CI(_15393_),
    .CO(_19374_),
    .S(_19375_));
 FA_X1 _40854_ (.A(_15477_),
    .B(_15458_),
    .CI(_15436_),
    .CO(_19376_),
    .S(_19377_));
 FA_X1 _40855_ (.A(_14820_),
    .B(_14797_),
    .CI(_14827_),
    .CO(_19378_),
    .S(_19379_));
 FA_X1 _40856_ (.A(_14849_),
    .B(_14856_),
    .CI(_14826_),
    .CO(_19380_),
    .S(_19381_));
 FA_X1 _40857_ (.A(_14877_),
    .B(_14883_),
    .CI(_14855_),
    .CO(_19382_),
    .S(_19383_));
 FA_X1 _40858_ (.A(_14908_),
    .B(_14901_),
    .CI(_14882_),
    .CO(_19384_),
    .S(_19385_));
 FA_X1 _40859_ (.A(_14921_),
    .B(_14926_),
    .CI(_14907_),
    .CO(_19386_),
    .S(_19387_));
 FA_X1 _40860_ (.A(_14935_),
    .B(_14943_),
    .CI(_14925_),
    .CO(_19388_),
    .S(_19389_));
 FA_X1 _40861_ (.A(_14948_),
    .B(_14956_),
    .CI(_14942_),
    .CO(_19390_),
    .S(_19391_));
 FA_X1 _40862_ (.A(_19392_),
    .B(_19393_),
    .CI(_14955_),
    .CO(_19394_),
    .S(_19395_));
 FA_X1 _40863_ (.A(_14967_),
    .B(_19396_),
    .CI(_14963_),
    .CO(\g_row[3].g_col[3].mult.stage1.dadda.t1[19] ),
    .S(\g_row[3].g_col[3].mult.stage1.dadda.t2[18] ));
 FA_X1 _40864_ (.A(_19397_),
    .B(_18850_),
    .CI(_19398_),
    .CO(_19399_),
    .S(_19400_));
 FA_X1 _40865_ (.A(_19401_),
    .B(_19402_),
    .CI(_19403_),
    .CO(_19404_),
    .S(_19405_));
 FA_X1 _40866_ (.A(_19406_),
    .B(_14708_),
    .CI(_19407_),
    .CO(\g_row[3].g_col[3].mult.stage1.dadda.t1[5] ),
    .S(\g_row[3].g_col[3].mult.stage1.dadda.t2[4] ));
 FA_X1 _40867_ (.A(_19408_),
    .B(_14718_),
    .CI(_19409_),
    .CO(_19410_),
    .S(_19411_));
 FA_X1 _40868_ (.A(_14717_),
    .B(_14723_),
    .CI(_19413_),
    .CO(_19414_),
    .S(_19415_));
 FA_X1 _40869_ (.A(_19416_),
    .B(_14749_),
    .CI(_19417_),
    .CO(_19418_),
    .S(_19419_));
 FA_X1 _40870_ (.A(_14764_),
    .B(_14773_),
    .CI(_14748_),
    .CO(_19420_),
    .S(_19421_));
 FA_X1 _40871_ (.A(_14792_),
    .B(_14798_),
    .CI(_14772_),
    .CO(_19422_),
    .S(_19423_));
 HA_X1 _40872_ (.A(_19424_),
    .B(_14210_),
    .CO(_19425_),
    .S(_19426_));
 HA_X1 _40873_ (.A(_14209_),
    .B(_14210_),
    .CO(_19427_),
    .S(_19428_));
 HA_X1 _40874_ (.A(_19429_),
    .B(_19430_),
    .CO(_19431_),
    .S(_19432_));
 HA_X1 _40875_ (.A(_19433_),
    .B(_19434_),
    .CO(_19435_),
    .S(_19436_));
 HA_X1 _40876_ (.A(_19437_),
    .B(_19438_),
    .CO(_19439_),
    .S(_19440_));
 HA_X1 _40877_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[0].g_col[0].mult.adder.b[20] ),
    .CO(_19441_),
    .S(_19442_));
 HA_X1 _40878_ (.A(\g_row[0].g_col[0].mult.adder.a[19] ),
    .B(\g_row[0].g_col[0].mult.adder.b[19] ),
    .CO(_19443_),
    .S(_19444_));
 HA_X1 _40879_ (.A(\g_row[0].g_col[0].mult.adder.a[18] ),
    .B(\g_row[0].g_col[0].mult.adder.b[18] ),
    .CO(_19445_),
    .S(_19446_));
 HA_X1 _40880_ (.A(\g_row[0].g_col[0].mult.adder.a[17] ),
    .B(\g_row[0].g_col[0].mult.adder.b[17] ),
    .CO(_19447_),
    .S(_19448_));
 HA_X1 _40881_ (.A(\g_row[0].g_col[0].mult.adder.a[16] ),
    .B(\g_row[0].g_col[0].mult.adder.b[16] ),
    .CO(_19449_),
    .S(_19450_));
 HA_X1 _40882_ (.A(\g_row[0].g_col[0].mult.adder.a[15] ),
    .B(\g_row[0].g_col[0].mult.adder.b[15] ),
    .CO(_19451_),
    .S(_19452_));
 HA_X1 _40883_ (.A(\g_row[0].g_col[0].mult.adder.a[14] ),
    .B(\g_row[0].g_col[0].mult.adder.b[14] ),
    .CO(_19453_),
    .S(_19454_));
 HA_X1 _40884_ (.A(\g_row[0].g_col[0].mult.adder.a[13] ),
    .B(\g_row[0].g_col[0].mult.adder.b[13] ),
    .CO(_19455_),
    .S(_19456_));
 HA_X1 _40885_ (.A(\g_row[0].g_col[0].mult.adder.a[12] ),
    .B(\g_row[0].g_col[0].mult.adder.b[12] ),
    .CO(_19457_),
    .S(_19458_));
 HA_X1 _40886_ (.A(\g_row[0].g_col[0].mult.adder.a[11] ),
    .B(\g_row[0].g_col[0].mult.adder.b[11] ),
    .CO(_19459_),
    .S(_19460_));
 HA_X1 _40887_ (.A(\g_row[0].g_col[0].mult.adder.a[10] ),
    .B(\g_row[0].g_col[0].mult.adder.b[10] ),
    .CO(_19461_),
    .S(_19462_));
 HA_X1 _40888_ (.A(\g_row[0].g_col[0].mult.adder.a[9] ),
    .B(\g_row[0].g_col[0].mult.adder.b[9] ),
    .CO(_19463_),
    .S(_19464_));
 HA_X1 _40889_ (.A(\g_row[0].g_col[0].mult.adder.a[8] ),
    .B(\g_row[0].g_col[0].mult.adder.b[8] ),
    .CO(_19465_),
    .S(_19466_));
 HA_X1 _40890_ (.A(\g_row[0].g_col[0].mult.adder.a[7] ),
    .B(\g_row[0].g_col[0].mult.adder.b[7] ),
    .CO(_19467_),
    .S(_19468_));
 HA_X1 _40891_ (.A(\g_row[0].g_col[0].mult.adder.a[6] ),
    .B(\g_row[0].g_col[0].mult.adder.b[6] ),
    .CO(_19469_),
    .S(_19470_));
 HA_X1 _40892_ (.A(\g_row[0].g_col[0].mult.adder.a[5] ),
    .B(\g_row[0].g_col[0].mult.adder.b[5] ),
    .CO(_19471_),
    .S(_19472_));
 HA_X1 _40893_ (.A(\g_row[0].g_col[0].mult.adder.a[4] ),
    .B(\g_row[0].g_col[0].mult.adder.b[4] ),
    .CO(_19473_),
    .S(_19474_));
 HA_X1 _40894_ (.A(\g_row[0].g_col[0].mult.adder.a[3] ),
    .B(\g_row[0].g_col[0].mult.adder.b[3] ),
    .CO(_19475_),
    .S(_19476_));
 HA_X1 _40895_ (.A(\g_row[0].g_col[0].mult.adder.a[2] ),
    .B(\g_row[0].g_col[0].mult.adder.b[2] ),
    .CO(_19477_),
    .S(_19478_));
 HA_X1 _40896_ (.A(\g_row[0].g_col[0].mult.adder.a[1] ),
    .B(\g_row[0].g_col[0].mult.adder.b[1] ),
    .CO(_19479_),
    .S(_19480_));
 HA_X1 _40897_ (.A(_19481_),
    .B(_19482_),
    .CO(_19483_),
    .S(_19484_));
 HA_X1 _40898_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19485_),
    .S(_19486_));
 HA_X1 _40899_ (.A(_19486_),
    .B(_19487_),
    .CO(_19488_),
    .S(_19489_));
 HA_X1 _40900_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19490_),
    .S(_19491_));
 HA_X1 _40901_ (.A(_19485_),
    .B(_19491_),
    .CO(_19492_),
    .S(_19493_));
 HA_X1 _40902_ (.A(_19494_),
    .B(_19495_),
    .CO(_19496_),
    .S(_19497_));
 HA_X1 _40903_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[0].g_col[1].mult.adder.b[20] ),
    .CO(_19498_),
    .S(_19499_));
 HA_X1 _40904_ (.A(\g_row[0].g_col[1].mult.adder.a[19] ),
    .B(\g_row[0].g_col[1].mult.adder.b[19] ),
    .CO(_19500_),
    .S(_19501_));
 HA_X1 _40905_ (.A(\g_row[0].g_col[1].mult.adder.a[18] ),
    .B(\g_row[0].g_col[1].mult.adder.b[18] ),
    .CO(_19502_),
    .S(_19503_));
 HA_X1 _40906_ (.A(\g_row[0].g_col[1].mult.adder.a[17] ),
    .B(\g_row[0].g_col[1].mult.adder.b[17] ),
    .CO(_19504_),
    .S(_19505_));
 HA_X1 _40907_ (.A(\g_row[0].g_col[1].mult.adder.a[16] ),
    .B(\g_row[0].g_col[1].mult.adder.b[16] ),
    .CO(_19506_),
    .S(_19507_));
 HA_X1 _40908_ (.A(\g_row[0].g_col[1].mult.adder.a[15] ),
    .B(\g_row[0].g_col[1].mult.adder.b[15] ),
    .CO(_19508_),
    .S(_19509_));
 HA_X1 _40909_ (.A(\g_row[0].g_col[1].mult.adder.a[14] ),
    .B(\g_row[0].g_col[1].mult.adder.b[14] ),
    .CO(_19510_),
    .S(_19511_));
 HA_X1 _40910_ (.A(\g_row[0].g_col[1].mult.adder.a[13] ),
    .B(\g_row[0].g_col[1].mult.adder.b[13] ),
    .CO(_19512_),
    .S(_19513_));
 HA_X1 _40911_ (.A(\g_row[0].g_col[1].mult.adder.a[12] ),
    .B(\g_row[0].g_col[1].mult.adder.b[12] ),
    .CO(_19514_),
    .S(_19515_));
 HA_X1 _40912_ (.A(\g_row[0].g_col[1].mult.adder.a[11] ),
    .B(\g_row[0].g_col[1].mult.adder.b[11] ),
    .CO(_19516_),
    .S(_19517_));
 HA_X1 _40913_ (.A(\g_row[0].g_col[1].mult.adder.a[10] ),
    .B(\g_row[0].g_col[1].mult.adder.b[10] ),
    .CO(_19518_),
    .S(_19519_));
 HA_X1 _40914_ (.A(\g_row[0].g_col[1].mult.adder.a[9] ),
    .B(\g_row[0].g_col[1].mult.adder.b[9] ),
    .CO(_19520_),
    .S(_19521_));
 HA_X1 _40915_ (.A(\g_row[0].g_col[1].mult.adder.a[8] ),
    .B(\g_row[0].g_col[1].mult.adder.b[8] ),
    .CO(_19522_),
    .S(_19523_));
 HA_X1 _40916_ (.A(\g_row[0].g_col[1].mult.adder.a[7] ),
    .B(\g_row[0].g_col[1].mult.adder.b[7] ),
    .CO(_19524_),
    .S(_19525_));
 HA_X1 _40917_ (.A(\g_row[0].g_col[1].mult.adder.a[6] ),
    .B(\g_row[0].g_col[1].mult.adder.b[6] ),
    .CO(_19526_),
    .S(_19527_));
 HA_X1 _40918_ (.A(\g_row[0].g_col[1].mult.adder.a[5] ),
    .B(\g_row[0].g_col[1].mult.adder.b[5] ),
    .CO(_19528_),
    .S(_19529_));
 HA_X1 _40919_ (.A(\g_row[0].g_col[1].mult.adder.a[4] ),
    .B(\g_row[0].g_col[1].mult.adder.b[4] ),
    .CO(_19530_),
    .S(_19531_));
 HA_X1 _40920_ (.A(\g_row[0].g_col[1].mult.adder.a[3] ),
    .B(\g_row[0].g_col[1].mult.adder.b[3] ),
    .CO(_19532_),
    .S(_19533_));
 HA_X1 _40921_ (.A(\g_row[0].g_col[1].mult.adder.a[2] ),
    .B(\g_row[0].g_col[1].mult.adder.b[2] ),
    .CO(_19534_),
    .S(_19535_));
 HA_X1 _40922_ (.A(\g_row[0].g_col[1].mult.adder.a[1] ),
    .B(\g_row[0].g_col[1].mult.adder.b[1] ),
    .CO(_19536_),
    .S(_19537_));
 HA_X1 _40923_ (.A(_19538_),
    .B(_19539_),
    .CO(_19540_),
    .S(_19541_));
 HA_X1 _40924_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19542_),
    .S(_19543_));
 HA_X1 _40925_ (.A(_19543_),
    .B(_19544_),
    .CO(_19545_),
    .S(_19546_));
 HA_X1 _40926_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19547_),
    .S(_19548_));
 HA_X1 _40927_ (.A(_19542_),
    .B(_19548_),
    .CO(_19549_),
    .S(_19550_));
 HA_X1 _40928_ (.A(_19551_),
    .B(_19552_),
    .CO(_19553_),
    .S(_19554_));
 HA_X1 _40929_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[0].g_col[2].mult.adder.b[20] ),
    .CO(_19555_),
    .S(_19556_));
 HA_X1 _40930_ (.A(\g_row[0].g_col[2].mult.adder.a[19] ),
    .B(\g_row[0].g_col[2].mult.adder.b[19] ),
    .CO(_19557_),
    .S(_19558_));
 HA_X1 _40931_ (.A(\g_row[0].g_col[2].mult.adder.a[18] ),
    .B(\g_row[0].g_col[2].mult.adder.b[18] ),
    .CO(_19559_),
    .S(_19560_));
 HA_X1 _40932_ (.A(\g_row[0].g_col[2].mult.adder.a[17] ),
    .B(\g_row[0].g_col[2].mult.adder.b[17] ),
    .CO(_19561_),
    .S(_19562_));
 HA_X1 _40933_ (.A(\g_row[0].g_col[2].mult.adder.a[16] ),
    .B(\g_row[0].g_col[2].mult.adder.b[16] ),
    .CO(_19563_),
    .S(_19564_));
 HA_X1 _40934_ (.A(\g_row[0].g_col[2].mult.adder.a[15] ),
    .B(\g_row[0].g_col[2].mult.adder.b[15] ),
    .CO(_19565_),
    .S(_19566_));
 HA_X1 _40935_ (.A(\g_row[0].g_col[2].mult.adder.a[14] ),
    .B(\g_row[0].g_col[2].mult.adder.b[14] ),
    .CO(_19567_),
    .S(_19568_));
 HA_X1 _40936_ (.A(\g_row[0].g_col[2].mult.adder.a[13] ),
    .B(\g_row[0].g_col[2].mult.adder.b[13] ),
    .CO(_19569_),
    .S(_19570_));
 HA_X1 _40937_ (.A(\g_row[0].g_col[2].mult.adder.a[12] ),
    .B(\g_row[0].g_col[2].mult.adder.b[12] ),
    .CO(_19571_),
    .S(_19572_));
 HA_X1 _40938_ (.A(\g_row[0].g_col[2].mult.adder.a[11] ),
    .B(\g_row[0].g_col[2].mult.adder.b[11] ),
    .CO(_19573_),
    .S(_19574_));
 HA_X1 _40939_ (.A(\g_row[0].g_col[2].mult.adder.a[10] ),
    .B(\g_row[0].g_col[2].mult.adder.b[10] ),
    .CO(_19575_),
    .S(_19576_));
 HA_X1 _40940_ (.A(\g_row[0].g_col[2].mult.adder.a[9] ),
    .B(\g_row[0].g_col[2].mult.adder.b[9] ),
    .CO(_19577_),
    .S(_19578_));
 HA_X1 _40941_ (.A(\g_row[0].g_col[2].mult.adder.a[8] ),
    .B(\g_row[0].g_col[2].mult.adder.b[8] ),
    .CO(_19579_),
    .S(_19580_));
 HA_X1 _40942_ (.A(\g_row[0].g_col[2].mult.adder.a[7] ),
    .B(\g_row[0].g_col[2].mult.adder.b[7] ),
    .CO(_19581_),
    .S(_19582_));
 HA_X1 _40943_ (.A(\g_row[0].g_col[2].mult.adder.a[6] ),
    .B(\g_row[0].g_col[2].mult.adder.b[6] ),
    .CO(_19583_),
    .S(_19584_));
 HA_X1 _40944_ (.A(\g_row[0].g_col[2].mult.adder.a[5] ),
    .B(\g_row[0].g_col[2].mult.adder.b[5] ),
    .CO(_19585_),
    .S(_19586_));
 HA_X1 _40945_ (.A(\g_row[0].g_col[2].mult.adder.a[4] ),
    .B(\g_row[0].g_col[2].mult.adder.b[4] ),
    .CO(_19587_),
    .S(_19588_));
 HA_X1 _40946_ (.A(\g_row[0].g_col[2].mult.adder.a[3] ),
    .B(\g_row[0].g_col[2].mult.adder.b[3] ),
    .CO(_19589_),
    .S(_19590_));
 HA_X1 _40947_ (.A(\g_row[0].g_col[2].mult.adder.a[2] ),
    .B(\g_row[0].g_col[2].mult.adder.b[2] ),
    .CO(_19591_),
    .S(_19592_));
 HA_X1 _40948_ (.A(\g_row[0].g_col[2].mult.adder.a[1] ),
    .B(\g_row[0].g_col[2].mult.adder.b[1] ),
    .CO(_19593_),
    .S(_19594_));
 HA_X1 _40949_ (.A(_19595_),
    .B(_19596_),
    .CO(_19597_),
    .S(_19598_));
 HA_X1 _40950_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19599_),
    .S(_19600_));
 HA_X1 _40951_ (.A(_19600_),
    .B(_19601_),
    .CO(_19602_),
    .S(_19603_));
 HA_X1 _40952_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19604_),
    .S(_19605_));
 HA_X1 _40953_ (.A(_19599_),
    .B(_19605_),
    .CO(_19606_),
    .S(_19607_));
 HA_X1 _40954_ (.A(_19608_),
    .B(_19609_),
    .CO(_19610_),
    .S(_19611_));
 HA_X1 _40955_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[0].g_col[3].mult.adder.b[20] ),
    .CO(_19612_),
    .S(_19613_));
 HA_X1 _40956_ (.A(\g_row[0].g_col[3].mult.adder.a[19] ),
    .B(\g_row[0].g_col[3].mult.adder.b[19] ),
    .CO(_19614_),
    .S(_19615_));
 HA_X1 _40957_ (.A(\g_row[0].g_col[3].mult.adder.a[18] ),
    .B(\g_row[0].g_col[3].mult.adder.b[18] ),
    .CO(_19616_),
    .S(_19617_));
 HA_X1 _40958_ (.A(\g_row[0].g_col[3].mult.adder.a[17] ),
    .B(\g_row[0].g_col[3].mult.adder.b[17] ),
    .CO(_19618_),
    .S(_19619_));
 HA_X1 _40959_ (.A(\g_row[0].g_col[3].mult.adder.a[16] ),
    .B(\g_row[0].g_col[3].mult.adder.b[16] ),
    .CO(_19620_),
    .S(_19621_));
 HA_X1 _40960_ (.A(\g_row[0].g_col[3].mult.adder.a[15] ),
    .B(\g_row[0].g_col[3].mult.adder.b[15] ),
    .CO(_19622_),
    .S(_19623_));
 HA_X1 _40961_ (.A(\g_row[0].g_col[3].mult.adder.a[14] ),
    .B(\g_row[0].g_col[3].mult.adder.b[14] ),
    .CO(_19624_),
    .S(_19625_));
 HA_X1 _40962_ (.A(\g_row[0].g_col[3].mult.adder.a[13] ),
    .B(\g_row[0].g_col[3].mult.adder.b[13] ),
    .CO(_19626_),
    .S(_19627_));
 HA_X1 _40963_ (.A(\g_row[0].g_col[3].mult.adder.a[12] ),
    .B(\g_row[0].g_col[3].mult.adder.b[12] ),
    .CO(_19628_),
    .S(_19629_));
 HA_X1 _40964_ (.A(\g_row[0].g_col[3].mult.adder.a[11] ),
    .B(\g_row[0].g_col[3].mult.adder.b[11] ),
    .CO(_19630_),
    .S(_19631_));
 HA_X1 _40965_ (.A(\g_row[0].g_col[3].mult.adder.a[10] ),
    .B(\g_row[0].g_col[3].mult.adder.b[10] ),
    .CO(_19632_),
    .S(_19633_));
 HA_X1 _40966_ (.A(\g_row[0].g_col[3].mult.adder.a[9] ),
    .B(\g_row[0].g_col[3].mult.adder.b[9] ),
    .CO(_19634_),
    .S(_19635_));
 HA_X1 _40967_ (.A(\g_row[0].g_col[3].mult.adder.a[8] ),
    .B(\g_row[0].g_col[3].mult.adder.b[8] ),
    .CO(_19636_),
    .S(_19637_));
 HA_X1 _40968_ (.A(\g_row[0].g_col[3].mult.adder.a[7] ),
    .B(\g_row[0].g_col[3].mult.adder.b[7] ),
    .CO(_19638_),
    .S(_19639_));
 HA_X1 _40969_ (.A(\g_row[0].g_col[3].mult.adder.a[6] ),
    .B(\g_row[0].g_col[3].mult.adder.b[6] ),
    .CO(_19640_),
    .S(_19641_));
 HA_X1 _40970_ (.A(\g_row[0].g_col[3].mult.adder.a[5] ),
    .B(\g_row[0].g_col[3].mult.adder.b[5] ),
    .CO(_19642_),
    .S(_19643_));
 HA_X1 _40971_ (.A(\g_row[0].g_col[3].mult.adder.a[4] ),
    .B(\g_row[0].g_col[3].mult.adder.b[4] ),
    .CO(_19644_),
    .S(_19645_));
 HA_X1 _40972_ (.A(\g_row[0].g_col[3].mult.adder.a[3] ),
    .B(\g_row[0].g_col[3].mult.adder.b[3] ),
    .CO(_19646_),
    .S(_19647_));
 HA_X1 _40973_ (.A(\g_row[0].g_col[3].mult.adder.a[2] ),
    .B(\g_row[0].g_col[3].mult.adder.b[2] ),
    .CO(_19648_),
    .S(_19649_));
 HA_X1 _40974_ (.A(\g_row[0].g_col[3].mult.adder.a[1] ),
    .B(\g_row[0].g_col[3].mult.adder.b[1] ),
    .CO(_19650_),
    .S(_19651_));
 HA_X1 _40975_ (.A(_19652_),
    .B(_19653_),
    .CO(_19654_),
    .S(_19655_));
 HA_X1 _40976_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19656_),
    .S(_19657_));
 HA_X1 _40977_ (.A(_19658_),
    .B(_19657_),
    .CO(_19659_),
    .S(_19660_));
 HA_X1 _40978_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19661_),
    .S(_19662_));
 HA_X1 _40979_ (.A(_19662_),
    .B(_19656_),
    .CO(_19663_),
    .S(_19664_));
 HA_X1 _40980_ (.A(_19665_),
    .B(_19666_),
    .CO(_19667_),
    .S(_19668_));
 HA_X1 _40981_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[1].g_col[0].mult.adder.b[20] ),
    .CO(_19669_),
    .S(_19670_));
 HA_X1 _40982_ (.A(\g_row[1].g_col[0].mult.adder.a[19] ),
    .B(\g_row[1].g_col[0].mult.adder.b[19] ),
    .CO(_19671_),
    .S(_19672_));
 HA_X1 _40983_ (.A(\g_row[1].g_col[0].mult.adder.a[18] ),
    .B(\g_row[1].g_col[0].mult.adder.b[18] ),
    .CO(_19673_),
    .S(_19674_));
 HA_X1 _40984_ (.A(\g_row[1].g_col[0].mult.adder.a[17] ),
    .B(\g_row[1].g_col[0].mult.adder.b[17] ),
    .CO(_19675_),
    .S(_19676_));
 HA_X1 _40985_ (.A(\g_row[1].g_col[0].mult.adder.a[16] ),
    .B(\g_row[1].g_col[0].mult.adder.b[16] ),
    .CO(_19677_),
    .S(_19678_));
 HA_X1 _40986_ (.A(\g_row[1].g_col[0].mult.adder.a[15] ),
    .B(\g_row[1].g_col[0].mult.adder.b[15] ),
    .CO(_19679_),
    .S(_19680_));
 HA_X1 _40987_ (.A(\g_row[1].g_col[0].mult.adder.a[14] ),
    .B(\g_row[1].g_col[0].mult.adder.b[14] ),
    .CO(_19681_),
    .S(_19682_));
 HA_X1 _40988_ (.A(\g_row[1].g_col[0].mult.adder.a[13] ),
    .B(\g_row[1].g_col[0].mult.adder.b[13] ),
    .CO(_19683_),
    .S(_19684_));
 HA_X1 _40989_ (.A(\g_row[1].g_col[0].mult.adder.a[12] ),
    .B(\g_row[1].g_col[0].mult.adder.b[12] ),
    .CO(_19685_),
    .S(_19686_));
 HA_X1 _40990_ (.A(\g_row[1].g_col[0].mult.adder.a[11] ),
    .B(\g_row[1].g_col[0].mult.adder.b[11] ),
    .CO(_19687_),
    .S(_19688_));
 HA_X1 _40991_ (.A(\g_row[1].g_col[0].mult.adder.a[10] ),
    .B(\g_row[1].g_col[0].mult.adder.b[10] ),
    .CO(_19689_),
    .S(_19690_));
 HA_X1 _40992_ (.A(\g_row[1].g_col[0].mult.adder.a[9] ),
    .B(\g_row[1].g_col[0].mult.adder.b[9] ),
    .CO(_19691_),
    .S(_19692_));
 HA_X1 _40993_ (.A(\g_row[1].g_col[0].mult.adder.a[8] ),
    .B(\g_row[1].g_col[0].mult.adder.b[8] ),
    .CO(_19693_),
    .S(_19694_));
 HA_X1 _40994_ (.A(\g_row[1].g_col[0].mult.adder.a[7] ),
    .B(\g_row[1].g_col[0].mult.adder.b[7] ),
    .CO(_19695_),
    .S(_19696_));
 HA_X1 _40995_ (.A(\g_row[1].g_col[0].mult.adder.a[6] ),
    .B(\g_row[1].g_col[0].mult.adder.b[6] ),
    .CO(_19697_),
    .S(_19698_));
 HA_X1 _40996_ (.A(\g_row[1].g_col[0].mult.adder.a[5] ),
    .B(\g_row[1].g_col[0].mult.adder.b[5] ),
    .CO(_19699_),
    .S(_19700_));
 HA_X1 _40997_ (.A(\g_row[1].g_col[0].mult.adder.a[4] ),
    .B(\g_row[1].g_col[0].mult.adder.b[4] ),
    .CO(_19701_),
    .S(_19702_));
 HA_X1 _40998_ (.A(\g_row[1].g_col[0].mult.adder.a[3] ),
    .B(\g_row[1].g_col[0].mult.adder.b[3] ),
    .CO(_19703_),
    .S(_19704_));
 HA_X1 _40999_ (.A(\g_row[1].g_col[0].mult.adder.a[2] ),
    .B(\g_row[1].g_col[0].mult.adder.b[2] ),
    .CO(_19705_),
    .S(_19706_));
 HA_X1 _41000_ (.A(\g_row[1].g_col[0].mult.adder.a[1] ),
    .B(\g_row[1].g_col[0].mult.adder.b[1] ),
    .CO(_19707_),
    .S(_19708_));
 HA_X1 _41001_ (.A(_19709_),
    .B(_19710_),
    .CO(_19711_),
    .S(_19712_));
 HA_X1 _41002_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[1].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19713_),
    .S(_19714_));
 HA_X1 _41003_ (.A(_19715_),
    .B(_19714_),
    .CO(_19716_),
    .S(_19717_));
 HA_X1 _41004_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[1].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19718_),
    .S(_19719_));
 HA_X1 _41005_ (.A(_19719_),
    .B(_19713_),
    .CO(_19720_),
    .S(_19721_));
 HA_X1 _41006_ (.A(_19722_),
    .B(_19723_),
    .CO(_19724_),
    .S(_19725_));
 HA_X1 _41007_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[1].g_col[1].mult.adder.b[20] ),
    .CO(_19726_),
    .S(_19727_));
 HA_X1 _41008_ (.A(\g_row[1].g_col[1].mult.adder.a[19] ),
    .B(\g_row[1].g_col[1].mult.adder.b[19] ),
    .CO(_19728_),
    .S(_19729_));
 HA_X1 _41009_ (.A(\g_row[1].g_col[1].mult.adder.a[18] ),
    .B(\g_row[1].g_col[1].mult.adder.b[18] ),
    .CO(_19730_),
    .S(_19731_));
 HA_X1 _41010_ (.A(\g_row[1].g_col[1].mult.adder.a[17] ),
    .B(\g_row[1].g_col[1].mult.adder.b[17] ),
    .CO(_19732_),
    .S(_19733_));
 HA_X1 _41011_ (.A(\g_row[1].g_col[1].mult.adder.a[16] ),
    .B(\g_row[1].g_col[1].mult.adder.b[16] ),
    .CO(_19734_),
    .S(_19735_));
 HA_X1 _41012_ (.A(\g_row[1].g_col[1].mult.adder.a[15] ),
    .B(\g_row[1].g_col[1].mult.adder.b[15] ),
    .CO(_19736_),
    .S(_19737_));
 HA_X1 _41013_ (.A(\g_row[1].g_col[1].mult.adder.a[14] ),
    .B(\g_row[1].g_col[1].mult.adder.b[14] ),
    .CO(_19738_),
    .S(_19739_));
 HA_X1 _41014_ (.A(\g_row[1].g_col[1].mult.adder.a[13] ),
    .B(\g_row[1].g_col[1].mult.adder.b[13] ),
    .CO(_19740_),
    .S(_19741_));
 HA_X1 _41015_ (.A(\g_row[1].g_col[1].mult.adder.a[12] ),
    .B(\g_row[1].g_col[1].mult.adder.b[12] ),
    .CO(_19742_),
    .S(_19743_));
 HA_X1 _41016_ (.A(\g_row[1].g_col[1].mult.adder.a[11] ),
    .B(\g_row[1].g_col[1].mult.adder.b[11] ),
    .CO(_19744_),
    .S(_19745_));
 HA_X1 _41017_ (.A(\g_row[1].g_col[1].mult.adder.a[10] ),
    .B(\g_row[1].g_col[1].mult.adder.b[10] ),
    .CO(_19746_),
    .S(_19747_));
 HA_X1 _41018_ (.A(\g_row[1].g_col[1].mult.adder.a[9] ),
    .B(\g_row[1].g_col[1].mult.adder.b[9] ),
    .CO(_19748_),
    .S(_19749_));
 HA_X1 _41019_ (.A(\g_row[1].g_col[1].mult.adder.a[8] ),
    .B(\g_row[1].g_col[1].mult.adder.b[8] ),
    .CO(_19750_),
    .S(_19751_));
 HA_X1 _41020_ (.A(\g_row[1].g_col[1].mult.adder.a[7] ),
    .B(\g_row[1].g_col[1].mult.adder.b[7] ),
    .CO(_19752_),
    .S(_19753_));
 HA_X1 _41021_ (.A(\g_row[1].g_col[1].mult.adder.a[6] ),
    .B(\g_row[1].g_col[1].mult.adder.b[6] ),
    .CO(_19754_),
    .S(_19755_));
 HA_X1 _41022_ (.A(\g_row[1].g_col[1].mult.adder.a[5] ),
    .B(\g_row[1].g_col[1].mult.adder.b[5] ),
    .CO(_19756_),
    .S(_19757_));
 HA_X1 _41023_ (.A(\g_row[1].g_col[1].mult.adder.a[4] ),
    .B(\g_row[1].g_col[1].mult.adder.b[4] ),
    .CO(_19758_),
    .S(_19759_));
 HA_X1 _41024_ (.A(\g_row[1].g_col[1].mult.adder.a[3] ),
    .B(\g_row[1].g_col[1].mult.adder.b[3] ),
    .CO(_19760_),
    .S(_19761_));
 HA_X1 _41025_ (.A(\g_row[1].g_col[1].mult.adder.a[2] ),
    .B(\g_row[1].g_col[1].mult.adder.b[2] ),
    .CO(_19762_),
    .S(_19763_));
 HA_X1 _41026_ (.A(\g_row[1].g_col[1].mult.adder.a[1] ),
    .B(\g_row[1].g_col[1].mult.adder.b[1] ),
    .CO(_19764_),
    .S(_19765_));
 HA_X1 _41027_ (.A(_19766_),
    .B(_19767_),
    .CO(_19768_),
    .S(_19769_));
 HA_X1 _41028_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[1].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19770_),
    .S(_19771_));
 HA_X1 _41029_ (.A(_19772_),
    .B(_19771_),
    .CO(_19773_),
    .S(_19774_));
 HA_X1 _41030_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[1].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19775_),
    .S(_19776_));
 HA_X1 _41031_ (.A(_19776_),
    .B(_19770_),
    .CO(_19777_),
    .S(_19778_));
 HA_X1 _41032_ (.A(_19779_),
    .B(_19780_),
    .CO(_19781_),
    .S(_19782_));
 HA_X1 _41033_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[1].g_col[2].mult.adder.b[20] ),
    .CO(_19783_),
    .S(_19784_));
 HA_X1 _41034_ (.A(\g_row[1].g_col[2].mult.adder.a[19] ),
    .B(\g_row[1].g_col[2].mult.adder.b[19] ),
    .CO(_19785_),
    .S(_19786_));
 HA_X1 _41035_ (.A(\g_row[1].g_col[2].mult.adder.a[18] ),
    .B(\g_row[1].g_col[2].mult.adder.b[18] ),
    .CO(_19787_),
    .S(_19788_));
 HA_X1 _41036_ (.A(\g_row[1].g_col[2].mult.adder.a[17] ),
    .B(\g_row[1].g_col[2].mult.adder.b[17] ),
    .CO(_19789_),
    .S(_19790_));
 HA_X1 _41037_ (.A(\g_row[1].g_col[2].mult.adder.a[16] ),
    .B(\g_row[1].g_col[2].mult.adder.b[16] ),
    .CO(_19791_),
    .S(_19792_));
 HA_X1 _41038_ (.A(\g_row[1].g_col[2].mult.adder.a[15] ),
    .B(\g_row[1].g_col[2].mult.adder.b[15] ),
    .CO(_19793_),
    .S(_19794_));
 HA_X1 _41039_ (.A(\g_row[1].g_col[2].mult.adder.a[14] ),
    .B(\g_row[1].g_col[2].mult.adder.b[14] ),
    .CO(_19795_),
    .S(_19796_));
 HA_X1 _41040_ (.A(\g_row[1].g_col[2].mult.adder.a[13] ),
    .B(\g_row[1].g_col[2].mult.adder.b[13] ),
    .CO(_19797_),
    .S(_19798_));
 HA_X1 _41041_ (.A(\g_row[1].g_col[2].mult.adder.a[12] ),
    .B(\g_row[1].g_col[2].mult.adder.b[12] ),
    .CO(_19799_),
    .S(_19800_));
 HA_X1 _41042_ (.A(\g_row[1].g_col[2].mult.adder.a[11] ),
    .B(\g_row[1].g_col[2].mult.adder.b[11] ),
    .CO(_19801_),
    .S(_19802_));
 HA_X1 _41043_ (.A(\g_row[1].g_col[2].mult.adder.a[10] ),
    .B(\g_row[1].g_col[2].mult.adder.b[10] ),
    .CO(_19803_),
    .S(_19804_));
 HA_X1 _41044_ (.A(\g_row[1].g_col[2].mult.adder.a[9] ),
    .B(\g_row[1].g_col[2].mult.adder.b[9] ),
    .CO(_19805_),
    .S(_19806_));
 HA_X1 _41045_ (.A(\g_row[1].g_col[2].mult.adder.a[8] ),
    .B(\g_row[1].g_col[2].mult.adder.b[8] ),
    .CO(_19807_),
    .S(_19808_));
 HA_X1 _41046_ (.A(\g_row[1].g_col[2].mult.adder.a[7] ),
    .B(\g_row[1].g_col[2].mult.adder.b[7] ),
    .CO(_19809_),
    .S(_19810_));
 HA_X1 _41047_ (.A(\g_row[1].g_col[2].mult.adder.a[6] ),
    .B(\g_row[1].g_col[2].mult.adder.b[6] ),
    .CO(_19811_),
    .S(_19812_));
 HA_X1 _41048_ (.A(\g_row[1].g_col[2].mult.adder.a[5] ),
    .B(\g_row[1].g_col[2].mult.adder.b[5] ),
    .CO(_19813_),
    .S(_19814_));
 HA_X1 _41049_ (.A(\g_row[1].g_col[2].mult.adder.a[4] ),
    .B(\g_row[1].g_col[2].mult.adder.b[4] ),
    .CO(_19815_),
    .S(_19816_));
 HA_X1 _41050_ (.A(\g_row[1].g_col[2].mult.adder.a[3] ),
    .B(\g_row[1].g_col[2].mult.adder.b[3] ),
    .CO(_19817_),
    .S(_19818_));
 HA_X1 _41051_ (.A(\g_row[1].g_col[2].mult.adder.a[2] ),
    .B(\g_row[1].g_col[2].mult.adder.b[2] ),
    .CO(_19819_),
    .S(_19820_));
 HA_X1 _41052_ (.A(\g_row[1].g_col[2].mult.adder.a[1] ),
    .B(\g_row[1].g_col[2].mult.adder.b[1] ),
    .CO(_19821_),
    .S(_19822_));
 HA_X1 _41053_ (.A(_19823_),
    .B(_19824_),
    .CO(_19825_),
    .S(_19826_));
 HA_X1 _41054_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[1].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19827_),
    .S(_19828_));
 HA_X1 _41055_ (.A(_19828_),
    .B(_19829_),
    .CO(_19830_),
    .S(_19831_));
 HA_X1 _41056_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[1].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19832_),
    .S(_19833_));
 HA_X1 _41057_ (.A(_19827_),
    .B(_19833_),
    .CO(_19834_),
    .S(_19835_));
 HA_X1 _41058_ (.A(_19836_),
    .B(_19837_),
    .CO(_19838_),
    .S(_19839_));
 HA_X1 _41059_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[1].g_col[3].mult.adder.b[20] ),
    .CO(_19840_),
    .S(_19841_));
 HA_X1 _41060_ (.A(\g_row[1].g_col[3].mult.adder.a[19] ),
    .B(\g_row[1].g_col[3].mult.adder.b[19] ),
    .CO(_19842_),
    .S(_19843_));
 HA_X1 _41061_ (.A(\g_row[1].g_col[3].mult.adder.a[18] ),
    .B(\g_row[1].g_col[3].mult.adder.b[18] ),
    .CO(_19844_),
    .S(_19845_));
 HA_X1 _41062_ (.A(\g_row[1].g_col[3].mult.adder.a[17] ),
    .B(\g_row[1].g_col[3].mult.adder.b[17] ),
    .CO(_19846_),
    .S(_19847_));
 HA_X1 _41063_ (.A(\g_row[1].g_col[3].mult.adder.a[16] ),
    .B(\g_row[1].g_col[3].mult.adder.b[16] ),
    .CO(_19848_),
    .S(_19849_));
 HA_X1 _41064_ (.A(\g_row[1].g_col[3].mult.adder.a[15] ),
    .B(\g_row[1].g_col[3].mult.adder.b[15] ),
    .CO(_19850_),
    .S(_19851_));
 HA_X1 _41065_ (.A(\g_row[1].g_col[3].mult.adder.a[14] ),
    .B(\g_row[1].g_col[3].mult.adder.b[14] ),
    .CO(_19852_),
    .S(_19853_));
 HA_X1 _41066_ (.A(\g_row[1].g_col[3].mult.adder.a[13] ),
    .B(\g_row[1].g_col[3].mult.adder.b[13] ),
    .CO(_19854_),
    .S(_19855_));
 HA_X1 _41067_ (.A(\g_row[1].g_col[3].mult.adder.a[12] ),
    .B(\g_row[1].g_col[3].mult.adder.b[12] ),
    .CO(_19856_),
    .S(_19857_));
 HA_X1 _41068_ (.A(\g_row[1].g_col[3].mult.adder.a[11] ),
    .B(\g_row[1].g_col[3].mult.adder.b[11] ),
    .CO(_19858_),
    .S(_19859_));
 HA_X1 _41069_ (.A(\g_row[1].g_col[3].mult.adder.a[10] ),
    .B(\g_row[1].g_col[3].mult.adder.b[10] ),
    .CO(_19860_),
    .S(_19861_));
 HA_X1 _41070_ (.A(\g_row[1].g_col[3].mult.adder.a[9] ),
    .B(\g_row[1].g_col[3].mult.adder.b[9] ),
    .CO(_19862_),
    .S(_19863_));
 HA_X1 _41071_ (.A(\g_row[1].g_col[3].mult.adder.a[8] ),
    .B(\g_row[1].g_col[3].mult.adder.b[8] ),
    .CO(_19864_),
    .S(_19865_));
 HA_X1 _41072_ (.A(\g_row[1].g_col[3].mult.adder.a[7] ),
    .B(\g_row[1].g_col[3].mult.adder.b[7] ),
    .CO(_19866_),
    .S(_19867_));
 HA_X1 _41073_ (.A(\g_row[1].g_col[3].mult.adder.a[6] ),
    .B(\g_row[1].g_col[3].mult.adder.b[6] ),
    .CO(_19868_),
    .S(_19869_));
 HA_X1 _41074_ (.A(\g_row[1].g_col[3].mult.adder.a[5] ),
    .B(\g_row[1].g_col[3].mult.adder.b[5] ),
    .CO(_19870_),
    .S(_19871_));
 HA_X1 _41075_ (.A(\g_row[1].g_col[3].mult.adder.a[4] ),
    .B(\g_row[1].g_col[3].mult.adder.b[4] ),
    .CO(_19872_),
    .S(_19873_));
 HA_X1 _41076_ (.A(\g_row[1].g_col[3].mult.adder.a[3] ),
    .B(\g_row[1].g_col[3].mult.adder.b[3] ),
    .CO(_19874_),
    .S(_19875_));
 HA_X1 _41077_ (.A(\g_row[1].g_col[3].mult.adder.a[2] ),
    .B(\g_row[1].g_col[3].mult.adder.b[2] ),
    .CO(_19876_),
    .S(_19877_));
 HA_X1 _41078_ (.A(\g_row[1].g_col[3].mult.adder.a[1] ),
    .B(\g_row[1].g_col[3].mult.adder.b[1] ),
    .CO(_19878_),
    .S(_19879_));
 HA_X1 _41079_ (.A(_19880_),
    .B(_19881_),
    .CO(_19882_),
    .S(_19883_));
 HA_X1 _41080_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[1].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19884_),
    .S(_19885_));
 HA_X1 _41081_ (.A(_19886_),
    .B(_19885_),
    .CO(_19887_),
    .S(_19888_));
 HA_X1 _41082_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[1].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19889_),
    .S(_19890_));
 HA_X1 _41083_ (.A(_19890_),
    .B(_19884_),
    .CO(_19891_),
    .S(_19892_));
 HA_X1 _41084_ (.A(_19893_),
    .B(_19894_),
    .CO(_19895_),
    .S(_19896_));
 HA_X1 _41085_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[2].g_col[0].mult.adder.b[20] ),
    .CO(_19897_),
    .S(_19898_));
 HA_X1 _41086_ (.A(\g_row[2].g_col[0].mult.adder.a[19] ),
    .B(\g_row[2].g_col[0].mult.adder.b[19] ),
    .CO(_19899_),
    .S(_19900_));
 HA_X1 _41087_ (.A(\g_row[2].g_col[0].mult.adder.a[18] ),
    .B(\g_row[2].g_col[0].mult.adder.b[18] ),
    .CO(_19901_),
    .S(_19902_));
 HA_X1 _41088_ (.A(\g_row[2].g_col[0].mult.adder.a[17] ),
    .B(\g_row[2].g_col[0].mult.adder.b[17] ),
    .CO(_19903_),
    .S(_19904_));
 HA_X1 _41089_ (.A(\g_row[2].g_col[0].mult.adder.a[16] ),
    .B(\g_row[2].g_col[0].mult.adder.b[16] ),
    .CO(_19905_),
    .S(_19906_));
 HA_X1 _41090_ (.A(\g_row[2].g_col[0].mult.adder.a[15] ),
    .B(\g_row[2].g_col[0].mult.adder.b[15] ),
    .CO(_19907_),
    .S(_19908_));
 HA_X1 _41091_ (.A(\g_row[2].g_col[0].mult.adder.a[14] ),
    .B(\g_row[2].g_col[0].mult.adder.b[14] ),
    .CO(_19909_),
    .S(_19910_));
 HA_X1 _41092_ (.A(\g_row[2].g_col[0].mult.adder.a[13] ),
    .B(\g_row[2].g_col[0].mult.adder.b[13] ),
    .CO(_19911_),
    .S(_19912_));
 HA_X1 _41093_ (.A(\g_row[2].g_col[0].mult.adder.a[12] ),
    .B(\g_row[2].g_col[0].mult.adder.b[12] ),
    .CO(_19913_),
    .S(_19914_));
 HA_X1 _41094_ (.A(\g_row[2].g_col[0].mult.adder.a[11] ),
    .B(\g_row[2].g_col[0].mult.adder.b[11] ),
    .CO(_19915_),
    .S(_19916_));
 HA_X1 _41095_ (.A(\g_row[2].g_col[0].mult.adder.a[10] ),
    .B(\g_row[2].g_col[0].mult.adder.b[10] ),
    .CO(_19917_),
    .S(_19918_));
 HA_X1 _41096_ (.A(\g_row[2].g_col[0].mult.adder.a[9] ),
    .B(\g_row[2].g_col[0].mult.adder.b[9] ),
    .CO(_19919_),
    .S(_19920_));
 HA_X1 _41097_ (.A(\g_row[2].g_col[0].mult.adder.a[8] ),
    .B(\g_row[2].g_col[0].mult.adder.b[8] ),
    .CO(_19921_),
    .S(_19922_));
 HA_X1 _41098_ (.A(\g_row[2].g_col[0].mult.adder.a[7] ),
    .B(\g_row[2].g_col[0].mult.adder.b[7] ),
    .CO(_19923_),
    .S(_19924_));
 HA_X1 _41099_ (.A(\g_row[2].g_col[0].mult.adder.a[6] ),
    .B(\g_row[2].g_col[0].mult.adder.b[6] ),
    .CO(_19925_),
    .S(_19926_));
 HA_X1 _41100_ (.A(\g_row[2].g_col[0].mult.adder.a[5] ),
    .B(\g_row[2].g_col[0].mult.adder.b[5] ),
    .CO(_19927_),
    .S(_19928_));
 HA_X1 _41101_ (.A(\g_row[2].g_col[0].mult.adder.a[4] ),
    .B(\g_row[2].g_col[0].mult.adder.b[4] ),
    .CO(_19929_),
    .S(_19930_));
 HA_X1 _41102_ (.A(\g_row[2].g_col[0].mult.adder.a[3] ),
    .B(\g_row[2].g_col[0].mult.adder.b[3] ),
    .CO(_19931_),
    .S(_19932_));
 HA_X1 _41103_ (.A(\g_row[2].g_col[0].mult.adder.a[2] ),
    .B(\g_row[2].g_col[0].mult.adder.b[2] ),
    .CO(_19933_),
    .S(_19934_));
 HA_X1 _41104_ (.A(\g_row[2].g_col[0].mult.adder.a[1] ),
    .B(\g_row[2].g_col[0].mult.adder.b[1] ),
    .CO(_19935_),
    .S(_19936_));
 HA_X1 _41105_ (.A(_19937_),
    .B(_19938_),
    .CO(_19939_),
    .S(_19940_));
 HA_X1 _41106_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[2].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19941_),
    .S(_19942_));
 HA_X1 _41107_ (.A(_19943_),
    .B(_19942_),
    .CO(_19944_),
    .S(_19945_));
 HA_X1 _41108_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[2].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_19946_),
    .S(_19947_));
 HA_X1 _41109_ (.A(_19947_),
    .B(_19941_),
    .CO(_19948_),
    .S(_19949_));
 HA_X1 _41110_ (.A(_19950_),
    .B(_19951_),
    .CO(_19952_),
    .S(_19953_));
 HA_X1 _41111_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[2].g_col[1].mult.adder.b[20] ),
    .CO(_19954_),
    .S(_19955_));
 HA_X1 _41112_ (.A(\g_row[2].g_col[1].mult.adder.a[19] ),
    .B(\g_row[2].g_col[1].mult.adder.b[19] ),
    .CO(_19956_),
    .S(_19957_));
 HA_X1 _41113_ (.A(\g_row[2].g_col[1].mult.adder.a[18] ),
    .B(\g_row[2].g_col[1].mult.adder.b[18] ),
    .CO(_19958_),
    .S(_19959_));
 HA_X1 _41114_ (.A(\g_row[2].g_col[1].mult.adder.a[17] ),
    .B(\g_row[2].g_col[1].mult.adder.b[17] ),
    .CO(_19960_),
    .S(_19961_));
 HA_X1 _41115_ (.A(\g_row[2].g_col[1].mult.adder.a[16] ),
    .B(\g_row[2].g_col[1].mult.adder.b[16] ),
    .CO(_19962_),
    .S(_19963_));
 HA_X1 _41116_ (.A(\g_row[2].g_col[1].mult.adder.a[15] ),
    .B(\g_row[2].g_col[1].mult.adder.b[15] ),
    .CO(_19964_),
    .S(_19965_));
 HA_X1 _41117_ (.A(\g_row[2].g_col[1].mult.adder.a[14] ),
    .B(\g_row[2].g_col[1].mult.adder.b[14] ),
    .CO(_19966_),
    .S(_19967_));
 HA_X1 _41118_ (.A(\g_row[2].g_col[1].mult.adder.a[13] ),
    .B(\g_row[2].g_col[1].mult.adder.b[13] ),
    .CO(_19968_),
    .S(_19969_));
 HA_X1 _41119_ (.A(\g_row[2].g_col[1].mult.adder.a[12] ),
    .B(\g_row[2].g_col[1].mult.adder.b[12] ),
    .CO(_19970_),
    .S(_19971_));
 HA_X1 _41120_ (.A(\g_row[2].g_col[1].mult.adder.a[11] ),
    .B(\g_row[2].g_col[1].mult.adder.b[11] ),
    .CO(_19972_),
    .S(_19973_));
 HA_X1 _41121_ (.A(\g_row[2].g_col[1].mult.adder.a[10] ),
    .B(\g_row[2].g_col[1].mult.adder.b[10] ),
    .CO(_19974_),
    .S(_19975_));
 HA_X1 _41122_ (.A(\g_row[2].g_col[1].mult.adder.a[9] ),
    .B(\g_row[2].g_col[1].mult.adder.b[9] ),
    .CO(_19976_),
    .S(_19977_));
 HA_X1 _41123_ (.A(\g_row[2].g_col[1].mult.adder.a[8] ),
    .B(\g_row[2].g_col[1].mult.adder.b[8] ),
    .CO(_19978_),
    .S(_19979_));
 HA_X1 _41124_ (.A(\g_row[2].g_col[1].mult.adder.a[7] ),
    .B(\g_row[2].g_col[1].mult.adder.b[7] ),
    .CO(_19980_),
    .S(_19981_));
 HA_X1 _41125_ (.A(\g_row[2].g_col[1].mult.adder.a[6] ),
    .B(\g_row[2].g_col[1].mult.adder.b[6] ),
    .CO(_19982_),
    .S(_19983_));
 HA_X1 _41126_ (.A(\g_row[2].g_col[1].mult.adder.a[5] ),
    .B(\g_row[2].g_col[1].mult.adder.b[5] ),
    .CO(_19984_),
    .S(_19985_));
 HA_X1 _41127_ (.A(\g_row[2].g_col[1].mult.adder.a[4] ),
    .B(\g_row[2].g_col[1].mult.adder.b[4] ),
    .CO(_19986_),
    .S(_19987_));
 HA_X1 _41128_ (.A(\g_row[2].g_col[1].mult.adder.a[3] ),
    .B(\g_row[2].g_col[1].mult.adder.b[3] ),
    .CO(_19988_),
    .S(_19989_));
 HA_X1 _41129_ (.A(\g_row[2].g_col[1].mult.adder.a[2] ),
    .B(\g_row[2].g_col[1].mult.adder.b[2] ),
    .CO(_19990_),
    .S(_19991_));
 HA_X1 _41130_ (.A(\g_row[2].g_col[1].mult.adder.a[1] ),
    .B(\g_row[2].g_col[1].mult.adder.b[1] ),
    .CO(_19992_),
    .S(_19993_));
 HA_X1 _41131_ (.A(_19994_),
    .B(_19995_),
    .CO(_19996_),
    .S(_19997_));
 HA_X1 _41132_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[2].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_19998_),
    .S(_19999_));
 HA_X1 _41133_ (.A(_19999_),
    .B(_20000_),
    .CO(_20001_),
    .S(_20002_));
 HA_X1 _41134_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[2].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20003_),
    .S(_20004_));
 HA_X1 _41135_ (.A(_20004_),
    .B(_19998_),
    .CO(_20005_),
    .S(_20006_));
 HA_X1 _41136_ (.A(_20007_),
    .B(_20008_),
    .CO(_20009_),
    .S(_20010_));
 HA_X1 _41137_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[2].g_col[2].mult.adder.b[20] ),
    .CO(_20011_),
    .S(_20012_));
 HA_X1 _41138_ (.A(\g_row[2].g_col[2].mult.adder.a[19] ),
    .B(\g_row[2].g_col[2].mult.adder.b[19] ),
    .CO(_20013_),
    .S(_20014_));
 HA_X1 _41139_ (.A(\g_row[2].g_col[2].mult.adder.a[18] ),
    .B(\g_row[2].g_col[2].mult.adder.b[18] ),
    .CO(_20015_),
    .S(_20016_));
 HA_X1 _41140_ (.A(\g_row[2].g_col[2].mult.adder.a[17] ),
    .B(\g_row[2].g_col[2].mult.adder.b[17] ),
    .CO(_20017_),
    .S(_20018_));
 HA_X1 _41141_ (.A(\g_row[2].g_col[2].mult.adder.a[16] ),
    .B(\g_row[2].g_col[2].mult.adder.b[16] ),
    .CO(_20019_),
    .S(_20020_));
 HA_X1 _41142_ (.A(\g_row[2].g_col[2].mult.adder.a[15] ),
    .B(\g_row[2].g_col[2].mult.adder.b[15] ),
    .CO(_20021_),
    .S(_20022_));
 HA_X1 _41143_ (.A(\g_row[2].g_col[2].mult.adder.a[14] ),
    .B(\g_row[2].g_col[2].mult.adder.b[14] ),
    .CO(_20023_),
    .S(_20024_));
 HA_X1 _41144_ (.A(\g_row[2].g_col[2].mult.adder.a[13] ),
    .B(\g_row[2].g_col[2].mult.adder.b[13] ),
    .CO(_20025_),
    .S(_20026_));
 HA_X1 _41145_ (.A(\g_row[2].g_col[2].mult.adder.a[12] ),
    .B(\g_row[2].g_col[2].mult.adder.b[12] ),
    .CO(_20027_),
    .S(_20028_));
 HA_X1 _41146_ (.A(\g_row[2].g_col[2].mult.adder.a[11] ),
    .B(\g_row[2].g_col[2].mult.adder.b[11] ),
    .CO(_20029_),
    .S(_20030_));
 HA_X1 _41147_ (.A(\g_row[2].g_col[2].mult.adder.a[10] ),
    .B(\g_row[2].g_col[2].mult.adder.b[10] ),
    .CO(_20031_),
    .S(_20032_));
 HA_X1 _41148_ (.A(\g_row[2].g_col[2].mult.adder.a[9] ),
    .B(\g_row[2].g_col[2].mult.adder.b[9] ),
    .CO(_20033_),
    .S(_20034_));
 HA_X1 _41149_ (.A(\g_row[2].g_col[2].mult.adder.a[8] ),
    .B(\g_row[2].g_col[2].mult.adder.b[8] ),
    .CO(_20035_),
    .S(_20036_));
 HA_X1 _41150_ (.A(\g_row[2].g_col[2].mult.adder.a[7] ),
    .B(\g_row[2].g_col[2].mult.adder.b[7] ),
    .CO(_20037_),
    .S(_20038_));
 HA_X1 _41151_ (.A(\g_row[2].g_col[2].mult.adder.a[6] ),
    .B(\g_row[2].g_col[2].mult.adder.b[6] ),
    .CO(_20039_),
    .S(_20040_));
 HA_X1 _41152_ (.A(\g_row[2].g_col[2].mult.adder.a[5] ),
    .B(\g_row[2].g_col[2].mult.adder.b[5] ),
    .CO(_20041_),
    .S(_20042_));
 HA_X1 _41153_ (.A(\g_row[2].g_col[2].mult.adder.a[4] ),
    .B(\g_row[2].g_col[2].mult.adder.b[4] ),
    .CO(_20043_),
    .S(_20044_));
 HA_X1 _41154_ (.A(\g_row[2].g_col[2].mult.adder.a[3] ),
    .B(\g_row[2].g_col[2].mult.adder.b[3] ),
    .CO(_20045_),
    .S(_20046_));
 HA_X1 _41155_ (.A(\g_row[2].g_col[2].mult.adder.a[2] ),
    .B(\g_row[2].g_col[2].mult.adder.b[2] ),
    .CO(_20047_),
    .S(_20048_));
 HA_X1 _41156_ (.A(\g_row[2].g_col[2].mult.adder.a[1] ),
    .B(\g_row[2].g_col[2].mult.adder.b[1] ),
    .CO(_20049_),
    .S(_20050_));
 HA_X1 _41157_ (.A(_20051_),
    .B(_20052_),
    .CO(_20053_),
    .S(_20054_));
 HA_X1 _41158_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[2].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20055_),
    .S(_20056_));
 HA_X1 _41159_ (.A(_20057_),
    .B(_20056_),
    .CO(_20058_),
    .S(_20059_));
 HA_X1 _41160_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[2].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20060_),
    .S(_20061_));
 HA_X1 _41161_ (.A(_20061_),
    .B(_20055_),
    .CO(_20062_),
    .S(_20063_));
 HA_X1 _41162_ (.A(_20064_),
    .B(_20065_),
    .CO(_20066_),
    .S(_20067_));
 HA_X1 _41163_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[2].g_col[3].mult.adder.b[20] ),
    .CO(_20068_),
    .S(_20069_));
 HA_X1 _41164_ (.A(\g_row[2].g_col[3].mult.adder.a[19] ),
    .B(\g_row[2].g_col[3].mult.adder.b[19] ),
    .CO(_20070_),
    .S(_20071_));
 HA_X1 _41165_ (.A(\g_row[2].g_col[3].mult.adder.a[18] ),
    .B(\g_row[2].g_col[3].mult.adder.b[18] ),
    .CO(_20072_),
    .S(_20073_));
 HA_X1 _41166_ (.A(\g_row[2].g_col[3].mult.adder.a[17] ),
    .B(\g_row[2].g_col[3].mult.adder.b[17] ),
    .CO(_20074_),
    .S(_20075_));
 HA_X1 _41167_ (.A(\g_row[2].g_col[3].mult.adder.a[16] ),
    .B(\g_row[2].g_col[3].mult.adder.b[16] ),
    .CO(_20076_),
    .S(_20077_));
 HA_X1 _41168_ (.A(\g_row[2].g_col[3].mult.adder.a[15] ),
    .B(\g_row[2].g_col[3].mult.adder.b[15] ),
    .CO(_20078_),
    .S(_20079_));
 HA_X1 _41169_ (.A(\g_row[2].g_col[3].mult.adder.a[14] ),
    .B(\g_row[2].g_col[3].mult.adder.b[14] ),
    .CO(_20080_),
    .S(_20081_));
 HA_X1 _41170_ (.A(\g_row[2].g_col[3].mult.adder.a[13] ),
    .B(\g_row[2].g_col[3].mult.adder.b[13] ),
    .CO(_20082_),
    .S(_20083_));
 HA_X1 _41171_ (.A(\g_row[2].g_col[3].mult.adder.a[12] ),
    .B(\g_row[2].g_col[3].mult.adder.b[12] ),
    .CO(_20084_),
    .S(_20085_));
 HA_X1 _41172_ (.A(\g_row[2].g_col[3].mult.adder.a[11] ),
    .B(\g_row[2].g_col[3].mult.adder.b[11] ),
    .CO(_20086_),
    .S(_20087_));
 HA_X1 _41173_ (.A(\g_row[2].g_col[3].mult.adder.a[10] ),
    .B(\g_row[2].g_col[3].mult.adder.b[10] ),
    .CO(_20088_),
    .S(_20089_));
 HA_X1 _41174_ (.A(\g_row[2].g_col[3].mult.adder.a[9] ),
    .B(\g_row[2].g_col[3].mult.adder.b[9] ),
    .CO(_20090_),
    .S(_20091_));
 HA_X1 _41175_ (.A(\g_row[2].g_col[3].mult.adder.a[8] ),
    .B(\g_row[2].g_col[3].mult.adder.b[8] ),
    .CO(_20092_),
    .S(_20093_));
 HA_X1 _41176_ (.A(\g_row[2].g_col[3].mult.adder.a[7] ),
    .B(\g_row[2].g_col[3].mult.adder.b[7] ),
    .CO(_20094_),
    .S(_20095_));
 HA_X1 _41177_ (.A(\g_row[2].g_col[3].mult.adder.a[6] ),
    .B(\g_row[2].g_col[3].mult.adder.b[6] ),
    .CO(_20096_),
    .S(_20097_));
 HA_X1 _41178_ (.A(\g_row[2].g_col[3].mult.adder.a[5] ),
    .B(\g_row[2].g_col[3].mult.adder.b[5] ),
    .CO(_20098_),
    .S(_20099_));
 HA_X1 _41179_ (.A(\g_row[2].g_col[3].mult.adder.a[4] ),
    .B(\g_row[2].g_col[3].mult.adder.b[4] ),
    .CO(_20100_),
    .S(_20101_));
 HA_X1 _41180_ (.A(\g_row[2].g_col[3].mult.adder.a[3] ),
    .B(\g_row[2].g_col[3].mult.adder.b[3] ),
    .CO(_20102_),
    .S(_20103_));
 HA_X1 _41181_ (.A(\g_row[2].g_col[3].mult.adder.a[2] ),
    .B(\g_row[2].g_col[3].mult.adder.b[2] ),
    .CO(_20104_),
    .S(_20105_));
 HA_X1 _41182_ (.A(\g_row[2].g_col[3].mult.adder.a[1] ),
    .B(\g_row[2].g_col[3].mult.adder.b[1] ),
    .CO(_20106_),
    .S(_20107_));
 HA_X1 _41183_ (.A(_20108_),
    .B(_20109_),
    .CO(_20110_),
    .S(_20111_));
 HA_X1 _41184_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[2].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20112_),
    .S(_20113_));
 HA_X1 _41185_ (.A(_20113_),
    .B(_20114_),
    .CO(_20115_),
    .S(_20116_));
 HA_X1 _41186_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[2].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20117_),
    .S(_20118_));
 HA_X1 _41187_ (.A(_20112_),
    .B(_20118_),
    .CO(_20119_),
    .S(_20120_));
 HA_X1 _41188_ (.A(_20121_),
    .B(_20122_),
    .CO(_20123_),
    .S(_20124_));
 HA_X1 _41189_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[3].g_col[0].mult.adder.b[20] ),
    .CO(_20125_),
    .S(_20126_));
 HA_X1 _41190_ (.A(\g_row[3].g_col[0].mult.adder.a[19] ),
    .B(\g_row[3].g_col[0].mult.adder.b[19] ),
    .CO(_20127_),
    .S(_20128_));
 HA_X1 _41191_ (.A(\g_row[3].g_col[0].mult.adder.a[18] ),
    .B(\g_row[3].g_col[0].mult.adder.b[18] ),
    .CO(_20129_),
    .S(_20130_));
 HA_X1 _41192_ (.A(\g_row[3].g_col[0].mult.adder.a[17] ),
    .B(\g_row[3].g_col[0].mult.adder.b[17] ),
    .CO(_20131_),
    .S(_20132_));
 HA_X1 _41193_ (.A(\g_row[3].g_col[0].mult.adder.a[16] ),
    .B(\g_row[3].g_col[0].mult.adder.b[16] ),
    .CO(_20133_),
    .S(_20134_));
 HA_X1 _41194_ (.A(\g_row[3].g_col[0].mult.adder.a[15] ),
    .B(\g_row[3].g_col[0].mult.adder.b[15] ),
    .CO(_20135_),
    .S(_20136_));
 HA_X1 _41195_ (.A(\g_row[3].g_col[0].mult.adder.a[14] ),
    .B(\g_row[3].g_col[0].mult.adder.b[14] ),
    .CO(_20137_),
    .S(_20138_));
 HA_X1 _41196_ (.A(\g_row[3].g_col[0].mult.adder.a[13] ),
    .B(\g_row[3].g_col[0].mult.adder.b[13] ),
    .CO(_20139_),
    .S(_20140_));
 HA_X1 _41197_ (.A(\g_row[3].g_col[0].mult.adder.a[12] ),
    .B(\g_row[3].g_col[0].mult.adder.b[12] ),
    .CO(_20141_),
    .S(_20142_));
 HA_X1 _41198_ (.A(\g_row[3].g_col[0].mult.adder.a[11] ),
    .B(\g_row[3].g_col[0].mult.adder.b[11] ),
    .CO(_20143_),
    .S(_20144_));
 HA_X1 _41199_ (.A(\g_row[3].g_col[0].mult.adder.a[10] ),
    .B(\g_row[3].g_col[0].mult.adder.b[10] ),
    .CO(_20145_),
    .S(_20146_));
 HA_X1 _41200_ (.A(\g_row[3].g_col[0].mult.adder.a[9] ),
    .B(\g_row[3].g_col[0].mult.adder.b[9] ),
    .CO(_20147_),
    .S(_20148_));
 HA_X1 _41201_ (.A(\g_row[3].g_col[0].mult.adder.a[8] ),
    .B(\g_row[3].g_col[0].mult.adder.b[8] ),
    .CO(_20149_),
    .S(_20150_));
 HA_X1 _41202_ (.A(\g_row[3].g_col[0].mult.adder.a[7] ),
    .B(\g_row[3].g_col[0].mult.adder.b[7] ),
    .CO(_20151_),
    .S(_20152_));
 HA_X1 _41203_ (.A(\g_row[3].g_col[0].mult.adder.a[6] ),
    .B(\g_row[3].g_col[0].mult.adder.b[6] ),
    .CO(_20153_),
    .S(_20154_));
 HA_X1 _41204_ (.A(\g_row[3].g_col[0].mult.adder.a[5] ),
    .B(\g_row[3].g_col[0].mult.adder.b[5] ),
    .CO(_20155_),
    .S(_20156_));
 HA_X1 _41205_ (.A(\g_row[3].g_col[0].mult.adder.a[4] ),
    .B(\g_row[3].g_col[0].mult.adder.b[4] ),
    .CO(_20157_),
    .S(_20158_));
 HA_X1 _41206_ (.A(\g_row[3].g_col[0].mult.adder.a[3] ),
    .B(\g_row[3].g_col[0].mult.adder.b[3] ),
    .CO(_20159_),
    .S(_20160_));
 HA_X1 _41207_ (.A(\g_row[3].g_col[0].mult.adder.a[2] ),
    .B(\g_row[3].g_col[0].mult.adder.b[2] ),
    .CO(_20161_),
    .S(_20162_));
 HA_X1 _41208_ (.A(\g_row[3].g_col[0].mult.adder.a[1] ),
    .B(\g_row[3].g_col[0].mult.adder.b[1] ),
    .CO(_20163_),
    .S(_20164_));
 HA_X1 _41209_ (.A(_20165_),
    .B(_20166_),
    .CO(_20167_),
    .S(_20168_));
 HA_X1 _41210_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[3].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20169_),
    .S(_20170_));
 HA_X1 _41211_ (.A(_20170_),
    .B(_20171_),
    .CO(_20172_),
    .S(_20173_));
 HA_X1 _41212_ (.A(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[3].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20174_),
    .S(_20175_));
 HA_X1 _41213_ (.A(_20175_),
    .B(_20169_),
    .CO(_20176_),
    .S(_20177_));
 HA_X1 _41214_ (.A(_20178_),
    .B(_20179_),
    .CO(_20180_),
    .S(_20181_));
 HA_X1 _41215_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[3].g_col[1].mult.adder.b[20] ),
    .CO(_20182_),
    .S(_20183_));
 HA_X1 _41216_ (.A(\g_row[3].g_col[1].mult.adder.a[19] ),
    .B(\g_row[3].g_col[1].mult.adder.b[19] ),
    .CO(_20184_),
    .S(_20185_));
 HA_X1 _41217_ (.A(\g_row[3].g_col[1].mult.adder.a[18] ),
    .B(\g_row[3].g_col[1].mult.adder.b[18] ),
    .CO(_20186_),
    .S(_20187_));
 HA_X1 _41218_ (.A(\g_row[3].g_col[1].mult.adder.a[17] ),
    .B(\g_row[3].g_col[1].mult.adder.b[17] ),
    .CO(_20188_),
    .S(_20189_));
 HA_X1 _41219_ (.A(\g_row[3].g_col[1].mult.adder.a[16] ),
    .B(\g_row[3].g_col[1].mult.adder.b[16] ),
    .CO(_20190_),
    .S(_20191_));
 HA_X1 _41220_ (.A(\g_row[3].g_col[1].mult.adder.a[15] ),
    .B(\g_row[3].g_col[1].mult.adder.b[15] ),
    .CO(_20192_),
    .S(_20193_));
 HA_X1 _41221_ (.A(\g_row[3].g_col[1].mult.adder.a[14] ),
    .B(\g_row[3].g_col[1].mult.adder.b[14] ),
    .CO(_20194_),
    .S(_20195_));
 HA_X1 _41222_ (.A(\g_row[3].g_col[1].mult.adder.a[13] ),
    .B(\g_row[3].g_col[1].mult.adder.b[13] ),
    .CO(_20196_),
    .S(_20197_));
 HA_X1 _41223_ (.A(\g_row[3].g_col[1].mult.adder.a[12] ),
    .B(\g_row[3].g_col[1].mult.adder.b[12] ),
    .CO(_20198_),
    .S(_20199_));
 HA_X1 _41224_ (.A(\g_row[3].g_col[1].mult.adder.a[11] ),
    .B(\g_row[3].g_col[1].mult.adder.b[11] ),
    .CO(_20200_),
    .S(_20201_));
 HA_X1 _41225_ (.A(\g_row[3].g_col[1].mult.adder.a[10] ),
    .B(\g_row[3].g_col[1].mult.adder.b[10] ),
    .CO(_20202_),
    .S(_20203_));
 HA_X1 _41226_ (.A(\g_row[3].g_col[1].mult.adder.a[9] ),
    .B(\g_row[3].g_col[1].mult.adder.b[9] ),
    .CO(_20204_),
    .S(_20205_));
 HA_X1 _41227_ (.A(\g_row[3].g_col[1].mult.adder.a[8] ),
    .B(\g_row[3].g_col[1].mult.adder.b[8] ),
    .CO(_20206_),
    .S(_20207_));
 HA_X1 _41228_ (.A(\g_row[3].g_col[1].mult.adder.a[7] ),
    .B(\g_row[3].g_col[1].mult.adder.b[7] ),
    .CO(_20208_),
    .S(_20209_));
 HA_X1 _41229_ (.A(\g_row[3].g_col[1].mult.adder.a[6] ),
    .B(\g_row[3].g_col[1].mult.adder.b[6] ),
    .CO(_20210_),
    .S(_20211_));
 HA_X1 _41230_ (.A(\g_row[3].g_col[1].mult.adder.a[5] ),
    .B(\g_row[3].g_col[1].mult.adder.b[5] ),
    .CO(_20212_),
    .S(_20213_));
 HA_X1 _41231_ (.A(\g_row[3].g_col[1].mult.adder.a[4] ),
    .B(\g_row[3].g_col[1].mult.adder.b[4] ),
    .CO(_20214_),
    .S(_20215_));
 HA_X1 _41232_ (.A(\g_row[3].g_col[1].mult.adder.a[3] ),
    .B(\g_row[3].g_col[1].mult.adder.b[3] ),
    .CO(_20216_),
    .S(_20217_));
 HA_X1 _41233_ (.A(\g_row[3].g_col[1].mult.adder.a[2] ),
    .B(\g_row[3].g_col[1].mult.adder.b[2] ),
    .CO(_20218_),
    .S(_20219_));
 HA_X1 _41234_ (.A(\g_row[3].g_col[1].mult.adder.a[1] ),
    .B(\g_row[3].g_col[1].mult.adder.b[1] ),
    .CO(_20220_),
    .S(_20221_));
 HA_X1 _41235_ (.A(_20222_),
    .B(_20223_),
    .CO(_20224_),
    .S(_20225_));
 HA_X1 _41236_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[3].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20226_),
    .S(_20227_));
 HA_X1 _41237_ (.A(_20228_),
    .B(_20227_),
    .CO(_20229_),
    .S(_20230_));
 HA_X1 _41238_ (.A(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[3].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20231_),
    .S(_20232_));
 HA_X1 _41239_ (.A(_20232_),
    .B(_20226_),
    .CO(_20233_),
    .S(_20234_));
 HA_X1 _41240_ (.A(_20235_),
    .B(_20236_),
    .CO(_20237_),
    .S(_20238_));
 HA_X1 _41241_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[3].g_col[2].mult.adder.b[20] ),
    .CO(_20239_),
    .S(_20240_));
 HA_X1 _41242_ (.A(\g_row[3].g_col[2].mult.adder.a[19] ),
    .B(\g_row[3].g_col[2].mult.adder.b[19] ),
    .CO(_20241_),
    .S(_20242_));
 HA_X1 _41243_ (.A(\g_row[3].g_col[2].mult.adder.a[18] ),
    .B(\g_row[3].g_col[2].mult.adder.b[18] ),
    .CO(_20243_),
    .S(_20244_));
 HA_X1 _41244_ (.A(\g_row[3].g_col[2].mult.adder.a[17] ),
    .B(\g_row[3].g_col[2].mult.adder.b[17] ),
    .CO(_20245_),
    .S(_20246_));
 HA_X1 _41245_ (.A(\g_row[3].g_col[2].mult.adder.a[16] ),
    .B(\g_row[3].g_col[2].mult.adder.b[16] ),
    .CO(_20247_),
    .S(_20248_));
 HA_X1 _41246_ (.A(\g_row[3].g_col[2].mult.adder.a[15] ),
    .B(\g_row[3].g_col[2].mult.adder.b[15] ),
    .CO(_20249_),
    .S(_20250_));
 HA_X1 _41247_ (.A(\g_row[3].g_col[2].mult.adder.a[14] ),
    .B(\g_row[3].g_col[2].mult.adder.b[14] ),
    .CO(_20251_),
    .S(_20252_));
 HA_X1 _41248_ (.A(\g_row[3].g_col[2].mult.adder.a[13] ),
    .B(\g_row[3].g_col[2].mult.adder.b[13] ),
    .CO(_20253_),
    .S(_20254_));
 HA_X1 _41249_ (.A(\g_row[3].g_col[2].mult.adder.a[12] ),
    .B(\g_row[3].g_col[2].mult.adder.b[12] ),
    .CO(_20255_),
    .S(_20256_));
 HA_X1 _41250_ (.A(\g_row[3].g_col[2].mult.adder.a[11] ),
    .B(\g_row[3].g_col[2].mult.adder.b[11] ),
    .CO(_20257_),
    .S(_20258_));
 HA_X1 _41251_ (.A(\g_row[3].g_col[2].mult.adder.a[10] ),
    .B(\g_row[3].g_col[2].mult.adder.b[10] ),
    .CO(_20259_),
    .S(_20260_));
 HA_X1 _41252_ (.A(\g_row[3].g_col[2].mult.adder.a[9] ),
    .B(\g_row[3].g_col[2].mult.adder.b[9] ),
    .CO(_20261_),
    .S(_20262_));
 HA_X1 _41253_ (.A(\g_row[3].g_col[2].mult.adder.a[8] ),
    .B(\g_row[3].g_col[2].mult.adder.b[8] ),
    .CO(_20263_),
    .S(_20264_));
 HA_X1 _41254_ (.A(\g_row[3].g_col[2].mult.adder.a[7] ),
    .B(\g_row[3].g_col[2].mult.adder.b[7] ),
    .CO(_20265_),
    .S(_20266_));
 HA_X1 _41255_ (.A(\g_row[3].g_col[2].mult.adder.a[6] ),
    .B(\g_row[3].g_col[2].mult.adder.b[6] ),
    .CO(_20267_),
    .S(_20268_));
 HA_X1 _41256_ (.A(\g_row[3].g_col[2].mult.adder.a[5] ),
    .B(\g_row[3].g_col[2].mult.adder.b[5] ),
    .CO(_20269_),
    .S(_20270_));
 HA_X1 _41257_ (.A(\g_row[3].g_col[2].mult.adder.a[4] ),
    .B(\g_row[3].g_col[2].mult.adder.b[4] ),
    .CO(_20271_),
    .S(_20272_));
 HA_X1 _41258_ (.A(\g_row[3].g_col[2].mult.adder.a[3] ),
    .B(\g_row[3].g_col[2].mult.adder.b[3] ),
    .CO(_20273_),
    .S(_20274_));
 HA_X1 _41259_ (.A(\g_row[3].g_col[2].mult.adder.a[2] ),
    .B(\g_row[3].g_col[2].mult.adder.b[2] ),
    .CO(_20275_),
    .S(_20276_));
 HA_X1 _41260_ (.A(\g_row[3].g_col[2].mult.adder.a[1] ),
    .B(\g_row[3].g_col[2].mult.adder.b[1] ),
    .CO(_20277_),
    .S(_20278_));
 HA_X1 _41261_ (.A(_20279_),
    .B(_20280_),
    .CO(_20281_),
    .S(_20282_));
 HA_X1 _41262_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[3].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20283_),
    .S(_20284_));
 HA_X1 _41263_ (.A(_20284_),
    .B(_20285_),
    .CO(_20286_),
    .S(_20287_));
 HA_X1 _41264_ (.A(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[3].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20288_),
    .S(_20289_));
 HA_X1 _41265_ (.A(_20283_),
    .B(_20289_),
    .CO(_20290_),
    .S(_20291_));
 HA_X1 _41266_ (.A(_20292_),
    .B(_20293_),
    .CO(_20294_),
    .S(_20295_));
 HA_X1 _41267_ (.A(\g_row[0].g_col[0].mult.adder.a[20] ),
    .B(\g_row[3].g_col[3].mult.adder.b[20] ),
    .CO(_20296_),
    .S(_20297_));
 HA_X1 _41268_ (.A(\g_row[3].g_col[3].mult.adder.a[19] ),
    .B(\g_row[3].g_col[3].mult.adder.b[19] ),
    .CO(_20298_),
    .S(_20299_));
 HA_X1 _41269_ (.A(\g_row[3].g_col[3].mult.adder.a[18] ),
    .B(\g_row[3].g_col[3].mult.adder.b[18] ),
    .CO(_20300_),
    .S(_20301_));
 HA_X1 _41270_ (.A(\g_row[3].g_col[3].mult.adder.a[17] ),
    .B(\g_row[3].g_col[3].mult.adder.b[17] ),
    .CO(_20302_),
    .S(_20303_));
 HA_X1 _41271_ (.A(\g_row[3].g_col[3].mult.adder.a[16] ),
    .B(\g_row[3].g_col[3].mult.adder.b[16] ),
    .CO(_20304_),
    .S(_20305_));
 HA_X1 _41272_ (.A(\g_row[3].g_col[3].mult.adder.a[15] ),
    .B(\g_row[3].g_col[3].mult.adder.b[15] ),
    .CO(_20306_),
    .S(_20307_));
 HA_X1 _41273_ (.A(\g_row[3].g_col[3].mult.adder.a[14] ),
    .B(\g_row[3].g_col[3].mult.adder.b[14] ),
    .CO(_20308_),
    .S(_20309_));
 HA_X1 _41274_ (.A(\g_row[3].g_col[3].mult.adder.a[13] ),
    .B(\g_row[3].g_col[3].mult.adder.b[13] ),
    .CO(_20310_),
    .S(_20311_));
 HA_X1 _41275_ (.A(\g_row[3].g_col[3].mult.adder.a[12] ),
    .B(\g_row[3].g_col[3].mult.adder.b[12] ),
    .CO(_20312_),
    .S(_20313_));
 HA_X1 _41276_ (.A(\g_row[3].g_col[3].mult.adder.a[11] ),
    .B(\g_row[3].g_col[3].mult.adder.b[11] ),
    .CO(_20314_),
    .S(_20315_));
 HA_X1 _41277_ (.A(\g_row[3].g_col[3].mult.adder.a[10] ),
    .B(\g_row[3].g_col[3].mult.adder.b[10] ),
    .CO(_20316_),
    .S(_20317_));
 HA_X1 _41278_ (.A(\g_row[3].g_col[3].mult.adder.a[9] ),
    .B(\g_row[3].g_col[3].mult.adder.b[9] ),
    .CO(_20318_),
    .S(_20319_));
 HA_X1 _41279_ (.A(\g_row[3].g_col[3].mult.adder.a[8] ),
    .B(\g_row[3].g_col[3].mult.adder.b[8] ),
    .CO(_20320_),
    .S(_20321_));
 HA_X1 _41280_ (.A(\g_row[3].g_col[3].mult.adder.a[7] ),
    .B(\g_row[3].g_col[3].mult.adder.b[7] ),
    .CO(_20322_),
    .S(_20323_));
 HA_X1 _41281_ (.A(\g_row[3].g_col[3].mult.adder.a[6] ),
    .B(\g_row[3].g_col[3].mult.adder.b[6] ),
    .CO(_20324_),
    .S(_20325_));
 HA_X1 _41282_ (.A(\g_row[3].g_col[3].mult.adder.a[5] ),
    .B(\g_row[3].g_col[3].mult.adder.b[5] ),
    .CO(_20326_),
    .S(_20327_));
 HA_X1 _41283_ (.A(\g_row[3].g_col[3].mult.adder.a[4] ),
    .B(\g_row[3].g_col[3].mult.adder.b[4] ),
    .CO(_20328_),
    .S(_20329_));
 HA_X1 _41284_ (.A(\g_row[3].g_col[3].mult.adder.a[3] ),
    .B(\g_row[3].g_col[3].mult.adder.b[3] ),
    .CO(_20330_),
    .S(_20331_));
 HA_X1 _41285_ (.A(\g_row[3].g_col[3].mult.adder.a[2] ),
    .B(\g_row[3].g_col[3].mult.adder.b[2] ),
    .CO(_20332_),
    .S(_20333_));
 HA_X1 _41286_ (.A(\g_row[3].g_col[3].mult.adder.a[1] ),
    .B(\g_row[3].g_col[3].mult.adder.b[1] ),
    .CO(_20334_),
    .S(_20335_));
 HA_X1 _41287_ (.A(_20336_),
    .B(_20337_),
    .CO(_20338_),
    .S(_20339_));
 HA_X1 _41288_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .B(\g_row[3].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .CO(_20340_),
    .S(_20341_));
 HA_X1 _41289_ (.A(_20341_),
    .B(_20342_),
    .CO(_20343_),
    .S(_20344_));
 HA_X1 _41290_ (.A(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .B(\g_row[3].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .CO(_20345_),
    .S(_20346_));
 HA_X1 _41291_ (.A(_20340_),
    .B(_20346_),
    .CO(_20347_),
    .S(_20348_));
 HA_X1 _41292_ (.A(_20349_),
    .B(_20350_),
    .CO(_20351_),
    .S(_20352_));
 HA_X1 _41293_ (.A(_20353_),
    .B(\g_reduce0[0].adder.a[13] ),
    .CO(_20354_),
    .S(_20355_));
 HA_X1 _41294_ (.A(_20356_),
    .B(\g_reduce0[0].adder.a[12] ),
    .CO(_20357_),
    .S(_20358_));
 HA_X1 _41295_ (.A(_20359_),
    .B(\g_reduce0[0].adder.a[11] ),
    .CO(_20360_),
    .S(_20361_));
 HA_X1 _41296_ (.A(_20362_),
    .B(\g_reduce0[0].adder.a[9] ),
    .CO(_20363_),
    .S(_20364_));
 HA_X1 _41297_ (.A(_20365_),
    .B(\g_reduce0[0].adder.a[8] ),
    .CO(_20366_),
    .S(_20367_));
 HA_X1 _41298_ (.A(_20368_),
    .B(\g_reduce0[0].adder.a[7] ),
    .CO(_20369_),
    .S(_20370_));
 HA_X1 _41299_ (.A(_20371_),
    .B(\g_reduce0[0].adder.a[6] ),
    .CO(_20372_),
    .S(_20373_));
 HA_X1 _41300_ (.A(_20374_),
    .B(\g_reduce0[0].adder.a[5] ),
    .CO(_20375_),
    .S(_20376_));
 HA_X1 _41301_ (.A(_20377_),
    .B(\g_reduce0[0].adder.a[4] ),
    .CO(_20378_),
    .S(_20379_));
 HA_X1 _41302_ (.A(_20380_),
    .B(\g_reduce0[0].adder.a[3] ),
    .CO(_20381_),
    .S(_20382_));
 HA_X1 _41303_ (.A(_20383_),
    .B(\g_reduce0[0].adder.a[2] ),
    .CO(_20384_),
    .S(_20385_));
 HA_X1 _41304_ (.A(_20386_),
    .B(\g_reduce0[0].adder.a[1] ),
    .CO(_20387_),
    .S(_20388_));
 HA_X1 _41305_ (.A(\g_reduce0[0].adder.b[0] ),
    .B(_20389_),
    .CO(_20390_),
    .S(_20391_));
 HA_X1 _41306_ (.A(\g_reduce0[0].adder.b[10] ),
    .B(_20392_),
    .CO(_20393_),
    .S(_20394_));
 HA_X1 _41307_ (.A(_20361_),
    .B(_20395_),
    .CO(_20396_),
    .S(_20397_));
 HA_X1 _41308_ (.A(_20398_),
    .B(\g_reduce0[0].adder.a[14] ),
    .CO(_20399_),
    .S(_20400_));
 HA_X1 _41309_ (.A(_14492_),
    .B(_14493_),
    .CO(_20401_),
    .S(_20402_));
 HA_X1 _41310_ (.A(_14493_),
    .B(_14497_),
    .CO(_20403_),
    .S(_20404_));
 HA_X1 _41311_ (.A(_20405_),
    .B(_20406_),
    .CO(_20407_),
    .S(_20408_));
 HA_X1 _41312_ (.A(_20409_),
    .B(_20410_),
    .CO(_20411_),
    .S(_20412_));
 HA_X1 _41313_ (.A(_20409_),
    .B(_20413_),
    .CO(_20414_),
    .S(_20415_));
 HA_X1 _41314_ (.A(_20416_),
    .B(_20417_),
    .CO(_20418_),
    .S(_20419_));
 HA_X1 _41315_ (.A(_20420_),
    .B(_20417_),
    .CO(_20421_),
    .S(_20422_));
 HA_X1 _41316_ (.A(_20423_),
    .B(_20424_),
    .CO(_20425_),
    .S(_20426_));
 HA_X1 _41317_ (.A(_20423_),
    .B(_20427_),
    .CO(_20428_),
    .S(_20429_));
 HA_X1 _41318_ (.A(_20430_),
    .B(_20431_),
    .CO(_20432_),
    .S(_20433_));
 HA_X1 _41319_ (.A(_20434_),
    .B(_20431_),
    .CO(_20435_),
    .S(_20436_));
 HA_X1 _41320_ (.A(_20437_),
    .B(_20438_),
    .CO(_20439_),
    .S(_20440_));
 HA_X1 _41321_ (.A(_20437_),
    .B(_20441_),
    .CO(_20442_),
    .S(_20443_));
 HA_X1 _41322_ (.A(_20444_),
    .B(_20445_),
    .CO(_20446_),
    .S(_20447_));
 HA_X1 _41323_ (.A(_20448_),
    .B(_20445_),
    .CO(_20449_),
    .S(_20450_));
 HA_X1 _41324_ (.A(_20406_),
    .B(_20451_),
    .CO(_20452_),
    .S(_20453_));
 HA_X1 _41325_ (.A(_20454_),
    .B(_20455_),
    .CO(_20456_),
    .S(_20457_));
 HA_X1 _41326_ (.A(_20458_),
    .B(_20455_),
    .CO(_20459_),
    .S(_20460_));
 HA_X1 _41327_ (.A(_20461_),
    .B(_20462_),
    .CO(_14491_),
    .S(_20463_));
 HA_X1 _41328_ (.A(_20462_),
    .B(_20464_),
    .CO(_14496_),
    .S(_20465_));
 HA_X1 _41329_ (.A(_20466_),
    .B(_20467_),
    .CO(_20468_),
    .S(_14506_));
 HA_X1 _41330_ (.A(_20466_),
    .B(_20469_),
    .CO(_20470_),
    .S(_20471_));
 HA_X1 _41331_ (.A(_20466_),
    .B(_20469_),
    .CO(_20472_),
    .S(_20473_));
 HA_X1 _41332_ (.A(_20474_),
    .B(_20475_),
    .CO(_20476_),
    .S(_20477_));
 HA_X1 _41333_ (.A(_20478_),
    .B(_20467_),
    .CO(_14502_),
    .S(_20479_));
 HA_X1 _41334_ (.A(_20480_),
    .B(_20481_),
    .CO(_20482_),
    .S(_20483_));
 HA_X1 _41335_ (.A(_20484_),
    .B(_14505_),
    .CO(_20485_),
    .S(_20486_));
 HA_X1 _41336_ (.A(_14505_),
    .B(_14506_),
    .CO(_20487_),
    .S(_20488_));
 HA_X1 _41337_ (.A(_20489_),
    .B(_20482_),
    .CO(_20490_),
    .S(_20491_));
 HA_X1 _41338_ (.A(_20492_),
    .B(_20493_),
    .CO(_20494_),
    .S(_20495_));
 HA_X1 _41339_ (.A(_20496_),
    .B(_20497_),
    .CO(_20498_),
    .S(_20499_));
 HA_X1 _41340_ (.A(\g_reduce0[10].adder.b[13] ),
    .B(_20500_),
    .CO(_20501_),
    .S(_20502_));
 HA_X1 _41341_ (.A(\g_reduce0[10].adder.b[12] ),
    .B(_20503_),
    .CO(_20504_),
    .S(_20505_));
 HA_X1 _41342_ (.A(\g_reduce0[10].adder.b[11] ),
    .B(_20506_),
    .CO(_20507_),
    .S(_20508_));
 HA_X1 _41343_ (.A(_20509_),
    .B(\g_reduce0[10].adder.a[10] ),
    .CO(_20510_),
    .S(_20511_));
 HA_X1 _41344_ (.A(\g_reduce0[10].adder.b[9] ),
    .B(_20512_),
    .CO(_20513_),
    .S(_20514_));
 HA_X1 _41345_ (.A(\g_reduce0[10].adder.b[8] ),
    .B(_20515_),
    .CO(_20516_),
    .S(_20517_));
 HA_X1 _41346_ (.A(\g_reduce0[10].adder.b[7] ),
    .B(_20518_),
    .CO(_20519_),
    .S(_20520_));
 HA_X1 _41347_ (.A(\g_reduce0[10].adder.b[6] ),
    .B(_20521_),
    .CO(_20522_),
    .S(_20523_));
 HA_X1 _41348_ (.A(\g_reduce0[10].adder.b[5] ),
    .B(_20524_),
    .CO(_20525_),
    .S(_20526_));
 HA_X1 _41349_ (.A(\g_reduce0[10].adder.b[4] ),
    .B(_20527_),
    .CO(_20528_),
    .S(_20529_));
 HA_X1 _41350_ (.A(\g_reduce0[10].adder.b[3] ),
    .B(_20530_),
    .CO(_20531_),
    .S(_20532_));
 HA_X1 _41351_ (.A(\g_reduce0[10].adder.b[2] ),
    .B(_20533_),
    .CO(_20534_),
    .S(_20535_));
 HA_X1 _41352_ (.A(\g_reduce0[10].adder.b[1] ),
    .B(_20536_),
    .CO(_20537_),
    .S(_20538_));
 HA_X1 _41353_ (.A(_20508_),
    .B(_20539_),
    .CO(_20540_),
    .S(_20541_));
 HA_X1 _41354_ (.A(\g_reduce0[10].adder.b[14] ),
    .B(_20542_),
    .CO(_20543_),
    .S(_20544_));
 HA_X1 _41355_ (.A(_14508_),
    .B(_14509_),
    .CO(_20545_),
    .S(_20546_));
 HA_X1 _41356_ (.A(_14512_),
    .B(_14509_),
    .CO(_20547_),
    .S(_20548_));
 HA_X1 _41357_ (.A(_20549_),
    .B(_20550_),
    .CO(_20551_),
    .S(_20552_));
 HA_X1 _41358_ (.A(_20553_),
    .B(_20554_),
    .CO(_20555_),
    .S(_20556_));
 HA_X1 _41359_ (.A(_20557_),
    .B(_20554_),
    .CO(_20558_),
    .S(_20559_));
 HA_X1 _41360_ (.A(_20560_),
    .B(_20561_),
    .CO(_20562_),
    .S(_20563_));
 HA_X1 _41361_ (.A(_20564_),
    .B(_20561_),
    .CO(_20565_),
    .S(_20566_));
 HA_X1 _41362_ (.A(_20567_),
    .B(_20568_),
    .CO(_20569_),
    .S(_20570_));
 HA_X1 _41363_ (.A(_20571_),
    .B(_20568_),
    .CO(_20572_),
    .S(_20573_));
 HA_X1 _41364_ (.A(_20574_),
    .B(_20575_),
    .CO(_20576_),
    .S(_20577_));
 HA_X1 _41365_ (.A(_20574_),
    .B(_20578_),
    .CO(_20579_),
    .S(_20580_));
 HA_X1 _41366_ (.A(_20581_),
    .B(_20582_),
    .CO(_20583_),
    .S(_20584_));
 HA_X1 _41367_ (.A(_20585_),
    .B(_20582_),
    .CO(_20586_),
    .S(_20587_));
 HA_X1 _41368_ (.A(_20588_),
    .B(_20589_),
    .CO(_20590_),
    .S(_20591_));
 HA_X1 _41369_ (.A(_20588_),
    .B(_20592_),
    .CO(_20593_),
    .S(_20594_));
 HA_X1 _41370_ (.A(_20549_),
    .B(_20595_),
    .CO(_20596_),
    .S(_20597_));
 HA_X1 _41371_ (.A(_20598_),
    .B(_20599_),
    .CO(_20600_),
    .S(_20601_));
 HA_X1 _41372_ (.A(_20598_),
    .B(_20602_),
    .CO(_20603_),
    .S(_20604_));
 HA_X1 _41373_ (.A(_20605_),
    .B(_20606_),
    .CO(_14507_),
    .S(_20607_));
 HA_X1 _41374_ (.A(_20606_),
    .B(_20608_),
    .CO(_14513_),
    .S(_20609_));
 HA_X1 _41375_ (.A(_20610_),
    .B(_20611_),
    .CO(_20612_),
    .S(_14517_));
 HA_X1 _41376_ (.A(_20610_),
    .B(_20613_),
    .CO(_20614_),
    .S(_20615_));
 HA_X1 _41377_ (.A(_20610_),
    .B(_20613_),
    .CO(_20616_),
    .S(_20617_));
 HA_X1 _41378_ (.A(_20618_),
    .B(_20619_),
    .CO(_20620_),
    .S(_20621_));
 HA_X1 _41379_ (.A(_20622_),
    .B(_20611_),
    .CO(_14521_),
    .S(_20623_));
 HA_X1 _41380_ (.A(_20624_),
    .B(_20625_),
    .CO(_20626_),
    .S(_20627_));
 HA_X1 _41381_ (.A(_20628_),
    .B(_14516_),
    .CO(_20629_),
    .S(_20630_));
 HA_X1 _41382_ (.A(_14516_),
    .B(_14517_),
    .CO(_20631_),
    .S(_20632_));
 HA_X1 _41383_ (.A(_20626_),
    .B(_20633_),
    .CO(_20634_),
    .S(_20635_));
 HA_X1 _41384_ (.A(_20636_),
    .B(_20637_),
    .CO(_20638_),
    .S(_20639_));
 HA_X1 _41385_ (.A(_20640_),
    .B(_20641_),
    .CO(_20642_),
    .S(_20643_));
 HA_X1 _41386_ (.A(_20644_),
    .B(_20645_),
    .CO(_14977_),
    .S(_20646_));
 HA_X1 _41387_ (.A(_20649_),
    .B(_20650_),
    .CO(_20647_),
    .S(_20651_));
 HA_X1 _41388_ (.A(_20652_),
    .B(_20653_),
    .CO(_20648_),
    .S(_14599_));
 HA_X1 _41389_ (.A(_20654_),
    .B(_20655_),
    .CO(_14600_),
    .S(_20656_));
 HA_X1 _41390_ (.A(net84),
    .B(net267),
    .CO(_14579_),
    .S(_20657_));
 HA_X1 _41391_ (.A(_20658_),
    .B(_20659_),
    .CO(_14621_),
    .S(_19087_));
 HA_X1 _41392_ (.A(_20661_),
    .B(_20662_),
    .CO(_20660_),
    .S(_19082_));
 HA_X1 _41393_ (.A(_20663_),
    .B(_20664_),
    .CO(_19081_),
    .S(_20665_));
 HA_X1 _41394_ (.A(_20666_),
    .B(_20667_),
    .CO(_19407_),
    .S(_20668_));
 HA_X1 _41395_ (.A(_20669_),
    .B(_20670_),
    .CO(_14674_),
    .S(_20671_));
 HA_X1 _41396_ (.A(_20673_),
    .B(_20674_),
    .CO(_20672_),
    .S(_20675_));
 HA_X1 _41397_ (.A(_20676_),
    .B(_20677_),
    .CO(_15143_),
    .S(_14673_));
 HA_X1 _41398_ (.A(_20678_),
    .B(_20679_),
    .CO(_20680_),
    .S(_19406_));
 HA_X1 _41399_ (.A(_20681_),
    .B(_20682_),
    .CO(_14729_),
    .S(_19412_));
 HA_X1 _41400_ (.A(_20683_),
    .B(_20684_),
    .CO(_14738_),
    .S(_20685_));
 HA_X1 _41401_ (.A(_20686_),
    .B(_20687_),
    .CO(_20688_),
    .S(_14737_));
 HA_X1 _41402_ (.A(_20689_),
    .B(_20690_),
    .CO(_14793_),
    .S(_20691_));
 HA_X1 _41403_ (.A(_20692_),
    .B(_20693_),
    .CO(_14803_),
    .S(_20694_));
 HA_X1 _41404_ (.A(_20695_),
    .B(_20696_),
    .CO(_14832_),
    .S(_14804_));
 HA_X1 _41405_ (.A(_20697_),
    .B(_20698_),
    .CO(_14866_),
    .S(_14833_));
 HA_X1 _41406_ (.A(net148),
    .B(net267),
    .CO(_14949_),
    .S(_20699_));
 HA_X1 _41407_ (.A(_20700_),
    .B(_20701_),
    .CO(_20702_),
    .S(_14978_));
 HA_X1 _41408_ (.A(_20704_),
    .B(_20705_),
    .CO(_14997_),
    .S(_20706_));
 HA_X1 _41409_ (.A(_20707_),
    .B(_20708_),
    .CO(_20709_),
    .S(_20710_));
 HA_X1 _41410_ (.A(_20711_),
    .B(_20712_),
    .CO(_20703_),
    .S(_20713_));
 HA_X1 _41411_ (.A(_20715_),
    .B(_20716_),
    .CO(_15081_),
    .S(_20717_));
 HA_X1 _41412_ (.A(_20718_),
    .B(_20719_),
    .CO(_15108_),
    .S(_15082_));
 HA_X1 _41413_ (.A(net36),
    .B(net275),
    .CO(_15165_),
    .S(_20720_));
 HA_X1 _41414_ (.A(_20721_),
    .B(_20722_),
    .CO(_15286_),
    .S(_20723_));
 HA_X1 _41415_ (.A(_20724_),
    .B(_20725_),
    .CO(_19218_),
    .S(_20726_));
 HA_X1 _41416_ (.A(_20727_),
    .B(_20728_),
    .CO(_19363_),
    .S(_20729_));
 HA_X1 _41417_ (.A(_20730_),
    .B(_20731_),
    .CO(_20732_),
    .S(_19362_));
 HA_X1 _41418_ (.A(_20733_),
    .B(_20734_),
    .CO(_15378_),
    .S(_20735_));
 HA_X1 _41419_ (.A(_20736_),
    .B(_20737_),
    .CO(_20738_),
    .S(_19219_));
 HA_X1 _41420_ (.A(_20739_),
    .B(_20740_),
    .CO(_20741_),
    .S(_20742_));
 HA_X1 _41421_ (.A(_20743_),
    .B(_20744_),
    .CO(_20745_),
    .S(_20746_));
 HA_X1 _41422_ (.A(_20747_),
    .B(_20748_),
    .CO(_15453_),
    .S(_20749_));
 HA_X1 _41423_ (.A(_20750_),
    .B(_20751_),
    .CO(_20752_),
    .S(_20753_));
 HA_X1 _41424_ (.A(_20754_),
    .B(_20755_),
    .CO(_15600_),
    .S(_20756_));
 HA_X1 _41425_ (.A(_20757_),
    .B(_20758_),
    .CO(_15533_),
    .S(_20759_));
 HA_X1 _41426_ (.A(_20760_),
    .B(_20761_),
    .CO(_15559_),
    .S(_15532_));
 HA_X1 _41427_ (.A(_20762_),
    .B(_20763_),
    .CO(_20714_),
    .S(_20764_));
 HA_X1 _41428_ (.A(net134),
    .B(net255),
    .CO(_15643_),
    .S(_20765_));
 HA_X1 _41429_ (.A(net68),
    .B(net255),
    .CO(_16477_),
    .S(_20766_));
 HA_X1 _41430_ (.A(_20767_),
    .B(_20768_),
    .CO(_19312_),
    .S(_20769_));
 HA_X1 _41431_ (.A(_20770_),
    .B(_20771_),
    .CO(_20772_),
    .S(_19313_));
 HA_X1 _41432_ (.A(_20773_),
    .B(_20774_),
    .CO(_15728_),
    .S(_19318_));
 HA_X1 _41433_ (.A(_20775_),
    .B(_20776_),
    .CO(_15750_),
    .S(_20777_));
 HA_X1 _41434_ (.A(_20778_),
    .B(_20779_),
    .CO(_20780_),
    .S(_15751_));
 HA_X1 _41435_ (.A(_20781_),
    .B(_20782_),
    .CO(_15795_),
    .S(_20783_));
 HA_X1 _41436_ (.A(_20784_),
    .B(_20785_),
    .CO(_15831_),
    .S(_20786_));
 HA_X1 _41437_ (.A(_20787_),
    .B(_20788_),
    .CO(_20789_),
    .S(_15832_));
 HA_X1 _41438_ (.A(_20790_),
    .B(_20791_),
    .CO(_15887_),
    .S(_20792_));
 HA_X1 _41439_ (.A(net117),
    .B(net243),
    .CO(_15970_),
    .S(_20793_));
 HA_X1 _41440_ (.A(_20794_),
    .B(_20795_),
    .CO(_16049_),
    .S(_16076_));
 HA_X1 _41441_ (.A(_20796_),
    .B(_20797_),
    .CO(_16077_),
    .S(_20798_));
 HA_X1 _41442_ (.A(_20800_),
    .B(_20801_),
    .CO(_20799_),
    .S(_20802_));
 HA_X1 _41443_ (.A(_20804_),
    .B(_20805_),
    .CO(_16147_),
    .S(_20806_));
 HA_X1 _41444_ (.A(_20807_),
    .B(_20808_),
    .CO(_20803_),
    .S(_16193_));
 HA_X1 _41445_ (.A(_20809_),
    .B(_20810_),
    .CO(_16194_),
    .S(_20811_));
 HA_X1 _41446_ (.A(_20813_),
    .B(_20814_),
    .CO(_16203_),
    .S(_20815_));
 HA_X1 _41447_ (.A(_20816_),
    .B(_20817_),
    .CO(_20812_),
    .S(_19129_));
 HA_X1 _41448_ (.A(_20818_),
    .B(_20819_),
    .CO(_19130_),
    .S(_19128_));
 HA_X1 _41449_ (.A(_20820_),
    .B(_20821_),
    .CO(_19263_),
    .S(_20822_));
 HA_X1 _41450_ (.A(_20823_),
    .B(_20824_),
    .CO(_20825_),
    .S(_19262_));
 HA_X1 _41451_ (.A(_20826_),
    .B(_20827_),
    .CO(_16249_),
    .S(_19268_));
 HA_X1 _41452_ (.A(_20828_),
    .B(_20829_),
    .CO(_16257_),
    .S(_20830_));
 HA_X1 _41453_ (.A(_20831_),
    .B(_20832_),
    .CO(_20833_),
    .S(_16258_));
 HA_X1 _41454_ (.A(_20834_),
    .B(_20835_),
    .CO(_20836_),
    .S(_20837_));
 HA_X1 _41455_ (.A(_20838_),
    .B(_20839_),
    .CO(_19175_),
    .S(_20840_));
 HA_X1 _41456_ (.A(_20841_),
    .B(_20842_),
    .CO(_16330_),
    .S(_20843_));
 HA_X1 _41457_ (.A(_20844_),
    .B(_20845_),
    .CO(_20846_),
    .S(_16329_));
 HA_X1 _41458_ (.A(_20847_),
    .B(_20848_),
    .CO(_16385_),
    .S(_20849_));
 HA_X1 _41459_ (.A(net101),
    .B(net275),
    .CO(_16465_),
    .S(_20850_));
 HA_X1 _41460_ (.A(net53),
    .B(net243),
    .CO(_16508_),
    .S(_20851_));
 HA_X1 _41461_ (.A(_20852_),
    .B(_20853_),
    .CO(_20854_),
    .S(_20855_));
 HA_X1 _41462_ (.A(_20856_),
    .B(_20857_),
    .CO(_20858_),
    .S(_20859_));
 HA_X1 _41463_ (.A(_20861_),
    .B(_20862_),
    .CO(_16543_),
    .S(_20863_));
 HA_X1 _41464_ (.A(_20864_),
    .B(_20865_),
    .CO(_20860_),
    .S(_19174_));
 HA_X1 _41465_ (.A(net221),
    .B(net275),
    .CO(_17640_),
    .S(_20866_));
 HA_X1 _41466_ (.A(_20867_),
    .B(_20868_),
    .CO(_16586_),
    .S(_20869_));
 HA_X1 _41467_ (.A(_20871_),
    .B(_20872_),
    .CO(_20870_),
    .S(_20873_));
 HA_X1 _41468_ (.A(_20876_),
    .B(_20877_),
    .CO(_16634_),
    .S(_20878_));
 HA_X1 _41469_ (.A(_20879_),
    .B(_20880_),
    .CO(_20874_),
    .S(_20881_));
 HA_X1 _41470_ (.A(_20882_),
    .B(_20883_),
    .CO(_20875_),
    .S(_18232_));
 HA_X1 _41471_ (.A(_20885_),
    .B(_20886_),
    .CO(_18590_),
    .S(_20887_));
 HA_X1 _41472_ (.A(_20888_),
    .B(_20889_),
    .CO(_16698_),
    .S(_20890_));
 HA_X1 _41473_ (.A(_20891_),
    .B(_20892_),
    .CO(_16766_),
    .S(_16812_));
 HA_X1 _41474_ (.A(_20893_),
    .B(_20894_),
    .CO(_16813_),
    .S(_20895_));
 HA_X1 _41475_ (.A(_20898_),
    .B(_20899_),
    .CO(_20897_),
    .S(_20900_));
 HA_X1 _41476_ (.A(_20902_),
    .B(_20903_),
    .CO(_18449_),
    .S(_20904_));
 HA_X1 _41477_ (.A(_20905_),
    .B(_20906_),
    .CO(_20901_),
    .S(_20907_));
 HA_X1 _41478_ (.A(_20908_),
    .B(_20909_),
    .CO(_18952_),
    .S(_18951_));
 HA_X1 _41479_ (.A(net204),
    .B(net275),
    .CO(_18249_),
    .S(_20910_));
 HA_X1 _41480_ (.A(_20911_),
    .B(_20912_),
    .CO(_16931_),
    .S(_20913_));
 HA_X1 _41481_ (.A(_20914_),
    .B(_20915_),
    .CO(_20916_),
    .S(_16932_));
 HA_X1 _41482_ (.A(_20918_),
    .B(_20919_),
    .CO(_16945_),
    .S(_20920_));
 HA_X1 _41483_ (.A(_20921_),
    .B(_20922_),
    .CO(_18381_),
    .S(_20923_));
 HA_X1 _41484_ (.A(_20924_),
    .B(_20925_),
    .CO(_17005_),
    .S(_17046_));
 HA_X1 _41485_ (.A(_20926_),
    .B(_20927_),
    .CO(_17047_),
    .S(_17585_));
 HA_X1 _41486_ (.A(_20928_),
    .B(_20929_),
    .CO(_17586_),
    .S(_20930_));
 HA_X1 _41487_ (.A(_20932_),
    .B(_20933_),
    .CO(_17078_),
    .S(_20934_));
 HA_X1 _41488_ (.A(_20935_),
    .B(_20936_),
    .CO(_20931_),
    .S(_18028_));
 HA_X1 _41489_ (.A(_20937_),
    .B(_20938_),
    .CO(_18545_),
    .S(_18863_));
 HA_X1 _41490_ (.A(_20940_),
    .B(_20941_),
    .CO(_17164_),
    .S(_20942_));
 HA_X1 _41491_ (.A(_20944_),
    .B(_20945_),
    .CO(_20943_),
    .S(_18013_));
 HA_X1 _41492_ (.A(_20946_),
    .B(_20947_),
    .CO(_18014_),
    .S(_20948_));
 HA_X1 _41493_ (.A(_20951_),
    .B(_20952_),
    .CO(_20949_),
    .S(_20953_));
 HA_X1 _41494_ (.A(_20954_),
    .B(_20955_),
    .CO(_20950_),
    .S(_17981_));
 HA_X1 _41495_ (.A(_20956_),
    .B(_20957_),
    .CO(_18496_),
    .S(_18818_));
 HA_X1 _41496_ (.A(_20960_),
    .B(_20961_),
    .CO(_17253_),
    .S(_20962_));
 HA_X1 _41497_ (.A(_20963_),
    .B(_20964_),
    .CO(_20965_),
    .S(_20966_));
 HA_X1 _41498_ (.A(_20967_),
    .B(_20968_),
    .CO(_20959_),
    .S(_17375_));
 HA_X1 _41499_ (.A(_20969_),
    .B(_20970_),
    .CO(_17329_),
    .S(_20971_));
 HA_X1 _41500_ (.A(_20972_),
    .B(_20973_),
    .CO(_17958_),
    .S(_17328_));
 HA_X1 _41501_ (.A(_20974_),
    .B(_20975_),
    .CO(_18765_),
    .S(_18763_));
 HA_X1 _41502_ (.A(_20976_),
    .B(_20977_),
    .CO(_17376_),
    .S(_20978_));
 HA_X1 _41503_ (.A(_20979_),
    .B(_20980_),
    .CO(_20981_),
    .S(_18994_));
 HA_X1 _41504_ (.A(_20983_),
    .B(_20984_),
    .CO(_18331_),
    .S(_20985_));
 HA_X1 _41505_ (.A(_20986_),
    .B(_20987_),
    .CO(_17479_),
    .S(_17460_));
 HA_X1 _41506_ (.A(_20988_),
    .B(_20989_),
    .CO(_17459_),
    .S(_20990_));
 HA_X1 _41507_ (.A(_20992_),
    .B(_20993_),
    .CO(_20991_),
    .S(_20994_));
 HA_X1 _41508_ (.A(_20995_),
    .B(_20996_),
    .CO(_20896_),
    .S(_20997_));
 HA_X1 _41509_ (.A(_20998_),
    .B(_20999_),
    .CO(_20917_),
    .S(_18380_));
 HA_X1 _41510_ (.A(_21001_),
    .B(_21002_),
    .CO(_18646_),
    .S(_21003_));
 HA_X1 _41511_ (.A(net21),
    .B(net267),
    .CO(_17680_),
    .S(_21004_));
 HA_X1 _41512_ (.A(_21005_),
    .B(_21006_),
    .CO(_17717_),
    .S(_17742_));
 HA_X1 _41513_ (.A(_21007_),
    .B(_21008_),
    .CO(_17741_),
    .S(_17763_));
 HA_X1 _41514_ (.A(_21009_),
    .B(_21010_),
    .CO(_17762_),
    .S(_21011_));
 HA_X1 _41515_ (.A(_21012_),
    .B(_21013_),
    .CO(_21014_),
    .S(_17802_));
 HA_X1 _41516_ (.A(_21015_),
    .B(_21016_),
    .CO(_17803_),
    .S(_21017_));
 HA_X1 _41517_ (.A(_21018_),
    .B(_21019_),
    .CO(_19036_),
    .S(_19033_));
 HA_X1 _41518_ (.A(net5),
    .B(net255),
    .CO(_18179_),
    .S(_21020_));
 HA_X1 _41519_ (.A(_21022_),
    .B(_21023_),
    .CO(_17888_),
    .S(_21024_));
 HA_X1 _41520_ (.A(_21025_),
    .B(_21026_),
    .CO(_21021_),
    .S(_21027_));
 HA_X1 _41521_ (.A(_21029_),
    .B(_21030_),
    .CO(_21028_),
    .S(_21031_));
 HA_X1 _41522_ (.A(_21032_),
    .B(_21033_),
    .CO(_18721_),
    .S(_18717_));
 HA_X1 _41523_ (.A(_21034_),
    .B(_21035_),
    .CO(_17982_),
    .S(_21036_));
 HA_X1 _41524_ (.A(net172),
    .B(net255),
    .CO(_17122_),
    .S(_21037_));
 HA_X1 _41525_ (.A(_21038_),
    .B(_21039_),
    .CO(_18029_),
    .S(_21040_));
 HA_X1 _41526_ (.A(_21041_),
    .B(_21042_),
    .CO(_21043_),
    .S(_18905_));
 HA_X1 _41527_ (.A(_21044_),
    .B(_21045_),
    .CO(_18091_),
    .S(_21046_));
 HA_X1 _41528_ (.A(_21048_),
    .B(_21049_),
    .CO(_18433_),
    .S(_21050_));
 HA_X1 _41529_ (.A(_21051_),
    .B(_21052_),
    .CO(_18201_),
    .S(_21053_));
 HA_X1 _41530_ (.A(_21054_),
    .B(_21055_),
    .CO(_18233_),
    .S(_21056_));
 HA_X1 _41531_ (.A(_21057_),
    .B(_21058_),
    .CO(_18812_),
    .S(_18811_));
 HA_X1 _41532_ (.A(_21059_),
    .B(_21060_),
    .CO(_18858_),
    .S(_18854_));
 HA_X1 _41533_ (.A(net187),
    .B(net267),
    .CO(_16986_),
    .S(_21061_));
 HA_X1 _41534_ (.A(net220),
    .B(net243),
    .CO(_16746_),
    .S(_21062_));
 HA_X1 _41535_ (.A(_21063_),
    .B(_21064_),
    .CO(_18995_),
    .S(_18991_));
 HA_X1 _41536_ (.A(_21065_),
    .B(_21066_),
    .CO(_18163_),
    .S(_21067_));
 HA_X1 _41537_ (.A(_21068_),
    .B(_21069_),
    .CO(_20982_),
    .S(_19037_));
 HA_X1 _41538_ (.A(_21070_),
    .B(_21071_),
    .CO(_18906_),
    .S(_18902_));
 HA_X1 _41539_ (.A(_21072_),
    .B(_21073_),
    .CO(_16963_),
    .S(_21074_));
 HA_X1 _41540_ (.A(_21075_),
    .B(_21076_),
    .CO(_21047_),
    .S(_18953_));
 HA_X1 _41541_ (.A(_21077_),
    .B(_21078_),
    .CO(_20958_),
    .S(_18813_));
 HA_X1 _41542_ (.A(_21079_),
    .B(_21080_),
    .CO(_20939_),
    .S(_18857_));
 HA_X1 _41543_ (.A(_21081_),
    .B(_21082_),
    .CO(_20884_),
    .S(_18720_));
 HA_X1 _41544_ (.A(_21083_),
    .B(_21084_),
    .CO(_21000_),
    .S(_18764_));
 HA_X1 _41545_ (.A(net149),
    .B(net243),
    .CO(_17359_),
    .S(_21085_));
 HA_X1 _41546_ (.A(_21086_),
    .B(_21087_),
    .CO(\g_row[0].g_col[0].mult.stage1.dadda.t1[3] ),
    .S(\g_row[0].g_col[0].mult.stage1.dadda.t2[2] ));
 HA_X1 _41547_ (.A(_21088_),
    .B(_21089_),
    .CO(\g_row[0].g_col[1].mult.stage1.dadda.t1[3] ),
    .S(\g_row[0].g_col[1].mult.stage1.dadda.t2[2] ));
 HA_X1 _41548_ (.A(_21090_),
    .B(_21091_),
    .CO(\g_row[0].g_col[2].mult.stage1.dadda.t1[3] ),
    .S(\g_row[0].g_col[2].mult.stage1.dadda.t2[2] ));
 HA_X1 _41549_ (.A(_21092_),
    .B(_21093_),
    .CO(\g_row[0].g_col[3].mult.stage1.dadda.t1[3] ),
    .S(\g_row[0].g_col[3].mult.stage1.dadda.t2[2] ));
 HA_X1 _41550_ (.A(_21094_),
    .B(_21095_),
    .CO(\g_row[1].g_col[0].mult.stage1.dadda.t1[3] ),
    .S(\g_row[1].g_col[0].mult.stage1.dadda.t2[2] ));
 HA_X1 _41551_ (.A(_21096_),
    .B(_21097_),
    .CO(\g_row[1].g_col[1].mult.stage1.dadda.t1[3] ),
    .S(\g_row[1].g_col[1].mult.stage1.dadda.t2[2] ));
 HA_X1 _41552_ (.A(_21098_),
    .B(_21099_),
    .CO(\g_row[1].g_col[2].mult.stage1.dadda.t1[3] ),
    .S(\g_row[1].g_col[2].mult.stage1.dadda.t2[2] ));
 HA_X1 _41553_ (.A(_21100_),
    .B(_21101_),
    .CO(\g_row[1].g_col[3].mult.stage1.dadda.t1[3] ),
    .S(\g_row[1].g_col[3].mult.stage1.dadda.t2[2] ));
 HA_X1 _41554_ (.A(_21102_),
    .B(_21103_),
    .CO(\g_row[2].g_col[0].mult.stage1.dadda.t1[3] ),
    .S(\g_row[2].g_col[0].mult.stage1.dadda.t2[2] ));
 HA_X1 _41555_ (.A(_21104_),
    .B(_21105_),
    .CO(\g_row[2].g_col[1].mult.stage1.dadda.t1[3] ),
    .S(\g_row[2].g_col[1].mult.stage1.dadda.t2[2] ));
 HA_X1 _41556_ (.A(_21106_),
    .B(_21107_),
    .CO(\g_row[2].g_col[2].mult.stage1.dadda.t1[3] ),
    .S(\g_row[2].g_col[2].mult.stage1.dadda.t2[2] ));
 HA_X1 _41557_ (.A(_21108_),
    .B(_21109_),
    .CO(\g_row[2].g_col[3].mult.stage1.dadda.t1[3] ),
    .S(\g_row[2].g_col[3].mult.stage1.dadda.t2[2] ));
 HA_X1 _41558_ (.A(_21110_),
    .B(_21111_),
    .CO(\g_row[3].g_col[0].mult.stage1.dadda.t1[3] ),
    .S(\g_row[3].g_col[0].mult.stage1.dadda.t2[2] ));
 HA_X1 _41559_ (.A(_21112_),
    .B(_21113_),
    .CO(\g_row[3].g_col[1].mult.stage1.dadda.t1[3] ),
    .S(\g_row[3].g_col[1].mult.stage1.dadda.t2[2] ));
 HA_X1 _41560_ (.A(_21114_),
    .B(_21115_),
    .CO(\g_row[3].g_col[2].mult.stage1.dadda.t1[3] ),
    .S(\g_row[3].g_col[2].mult.stage1.dadda.t2[2] ));
 HA_X1 _41561_ (.A(_21116_),
    .B(_21117_),
    .CO(\g_row[3].g_col[3].mult.stage1.dadda.t1[3] ),
    .S(\g_row[3].g_col[3].mult.stage1.dadda.t2[2] ));
 HA_X1 _41562_ (.A(\g_reduce0[12].adder.b[13] ),
    .B(_21118_),
    .CO(_21119_),
    .S(_21120_));
 HA_X1 _41563_ (.A(\g_reduce0[12].adder.b[12] ),
    .B(_21121_),
    .CO(_21122_),
    .S(_21123_));
 HA_X1 _41564_ (.A(\g_reduce0[12].adder.b[11] ),
    .B(_21124_),
    .CO(_21125_),
    .S(_21126_));
 HA_X1 _41565_ (.A(_21127_),
    .B(\g_reduce0[12].adder.a[10] ),
    .CO(_21128_),
    .S(_21129_));
 HA_X1 _41566_ (.A(\g_reduce0[12].adder.b[9] ),
    .B(_21130_),
    .CO(_21131_),
    .S(_21132_));
 HA_X1 _41567_ (.A(\g_reduce0[12].adder.b[8] ),
    .B(_21133_),
    .CO(_21134_),
    .S(_21135_));
 HA_X1 _41568_ (.A(\g_reduce0[12].adder.b[7] ),
    .B(_21136_),
    .CO(_21137_),
    .S(_21138_));
 HA_X1 _41569_ (.A(\g_reduce0[12].adder.b[6] ),
    .B(_21139_),
    .CO(_21140_),
    .S(_21141_));
 HA_X1 _41570_ (.A(\g_reduce0[12].adder.b[5] ),
    .B(_21142_),
    .CO(_21143_),
    .S(_21144_));
 HA_X1 _41571_ (.A(\g_reduce0[12].adder.b[4] ),
    .B(_21145_),
    .CO(_21146_),
    .S(_21147_));
 HA_X1 _41572_ (.A(\g_reduce0[12].adder.b[3] ),
    .B(_21148_),
    .CO(_21149_),
    .S(_21150_));
 HA_X1 _41573_ (.A(\g_reduce0[12].adder.b[2] ),
    .B(_21151_),
    .CO(_21152_),
    .S(_21153_));
 HA_X1 _41574_ (.A(\g_reduce0[12].adder.b[1] ),
    .B(_21154_),
    .CO(_21155_),
    .S(_21156_));
 HA_X1 _41575_ (.A(_21157_),
    .B(_21126_),
    .CO(_21158_),
    .S(_21159_));
 HA_X1 _41576_ (.A(\g_reduce0[12].adder.b[14] ),
    .B(_21160_),
    .CO(_21161_),
    .S(_21162_));
 HA_X1 _41577_ (.A(_14059_),
    .B(_14060_),
    .CO(_21163_),
    .S(_21164_));
 HA_X1 _41578_ (.A(_14060_),
    .B(_14064_),
    .CO(_21165_),
    .S(_21166_));
 HA_X1 _41579_ (.A(_21167_),
    .B(_21168_),
    .CO(_21169_),
    .S(_21170_));
 HA_X1 _41580_ (.A(_21171_),
    .B(_21172_),
    .CO(_21173_),
    .S(_21174_));
 HA_X1 _41581_ (.A(_21171_),
    .B(_21175_),
    .CO(_21176_),
    .S(_21177_));
 HA_X1 _41582_ (.A(_21178_),
    .B(_21179_),
    .CO(_21180_),
    .S(_21181_));
 HA_X1 _41583_ (.A(_21182_),
    .B(_21179_),
    .CO(_21183_),
    .S(_21184_));
 HA_X1 _41584_ (.A(_21185_),
    .B(_21186_),
    .CO(_21187_),
    .S(_21188_));
 HA_X1 _41585_ (.A(_21189_),
    .B(_21186_),
    .CO(_21190_),
    .S(_21191_));
 HA_X1 _41586_ (.A(_21192_),
    .B(_21193_),
    .CO(_21194_),
    .S(_21195_));
 HA_X1 _41587_ (.A(_21192_),
    .B(_21196_),
    .CO(_21197_),
    .S(_21198_));
 HA_X1 _41588_ (.A(_21199_),
    .B(_21200_),
    .CO(_21201_),
    .S(_21202_));
 HA_X1 _41589_ (.A(_21199_),
    .B(_21203_),
    .CO(_21204_),
    .S(_21205_));
 HA_X1 _41590_ (.A(_21206_),
    .B(_21207_),
    .CO(_21208_),
    .S(_21209_));
 HA_X1 _41591_ (.A(_21210_),
    .B(_21207_),
    .CO(_21211_),
    .S(_21212_));
 HA_X1 _41592_ (.A(_21213_),
    .B(_21167_),
    .CO(_21214_),
    .S(_21215_));
 HA_X1 _41593_ (.A(_21216_),
    .B(_21217_),
    .CO(_21218_),
    .S(_21219_));
 HA_X1 _41594_ (.A(_21216_),
    .B(_21220_),
    .CO(_21221_),
    .S(_21222_));
 HA_X1 _41595_ (.A(_21223_),
    .B(_21224_),
    .CO(_14058_),
    .S(_21225_));
 HA_X1 _41596_ (.A(_21224_),
    .B(_21226_),
    .CO(_14063_),
    .S(_21227_));
 HA_X1 _41597_ (.A(_21228_),
    .B(_21229_),
    .CO(_21230_),
    .S(_14068_));
 HA_X1 _41598_ (.A(_21228_),
    .B(_21231_),
    .CO(_21232_),
    .S(_21233_));
 HA_X1 _41599_ (.A(_21228_),
    .B(_21231_),
    .CO(_21234_),
    .S(_21235_));
 HA_X1 _41600_ (.A(_21236_),
    .B(_21237_),
    .CO(_21238_),
    .S(_21239_));
 HA_X1 _41601_ (.A(_21240_),
    .B(_21229_),
    .CO(_14072_),
    .S(_21241_));
 HA_X1 _41602_ (.A(_21242_),
    .B(_21243_),
    .CO(_21244_),
    .S(_21245_));
 HA_X1 _41603_ (.A(_14067_),
    .B(_21246_),
    .CO(_21247_),
    .S(_21248_));
 HA_X1 _41604_ (.A(_14067_),
    .B(_14068_),
    .CO(_21249_),
    .S(_21250_));
 HA_X1 _41605_ (.A(_21251_),
    .B(_21244_),
    .CO(_21252_),
    .S(_21253_));
 HA_X1 _41606_ (.A(_21254_),
    .B(_21255_),
    .CO(_21256_),
    .S(_21257_));
 HA_X1 _41607_ (.A(_21258_),
    .B(_21259_),
    .CO(_21260_),
    .S(_21261_));
 HA_X1 _41608_ (.A(_21262_),
    .B(\g_reduce0[14].adder.a[13] ),
    .CO(_21263_),
    .S(_21264_));
 HA_X1 _41609_ (.A(_21265_),
    .B(\g_reduce0[14].adder.a[12] ),
    .CO(_21266_),
    .S(_21267_));
 HA_X1 _41610_ (.A(_21268_),
    .B(\g_reduce0[14].adder.a[11] ),
    .CO(_21269_),
    .S(_21270_));
 HA_X1 _41611_ (.A(_21271_),
    .B(\g_reduce0[14].adder.a[9] ),
    .CO(_21272_),
    .S(_21273_));
 HA_X1 _41612_ (.A(_21274_),
    .B(\g_reduce0[14].adder.a[8] ),
    .CO(_21275_),
    .S(_21276_));
 HA_X1 _41613_ (.A(_21277_),
    .B(\g_reduce0[14].adder.a[7] ),
    .CO(_21278_),
    .S(_21279_));
 HA_X1 _41614_ (.A(_21280_),
    .B(\g_reduce0[14].adder.a[6] ),
    .CO(_21281_),
    .S(_21282_));
 HA_X1 _41615_ (.A(_21283_),
    .B(\g_reduce0[14].adder.a[5] ),
    .CO(_21284_),
    .S(_21285_));
 HA_X1 _41616_ (.A(_21286_),
    .B(\g_reduce0[14].adder.a[4] ),
    .CO(_21287_),
    .S(_21288_));
 HA_X1 _41617_ (.A(_21289_),
    .B(\g_reduce0[14].adder.a[3] ),
    .CO(_21290_),
    .S(_21291_));
 HA_X1 _41618_ (.A(_21292_),
    .B(\g_reduce0[14].adder.a[2] ),
    .CO(_21293_),
    .S(_21294_));
 HA_X1 _41619_ (.A(_21295_),
    .B(\g_reduce0[14].adder.a[1] ),
    .CO(_21296_),
    .S(_21297_));
 HA_X1 _41620_ (.A(\g_reduce0[14].adder.b[0] ),
    .B(_21298_),
    .CO(_21299_),
    .S(_21300_));
 HA_X1 _41621_ (.A(\g_reduce0[14].adder.b[10] ),
    .B(_21301_),
    .CO(_21302_),
    .S(_21303_));
 HA_X1 _41622_ (.A(_21270_),
    .B(_21304_),
    .CO(_21305_),
    .S(_21306_));
 HA_X1 _41623_ (.A(_21307_),
    .B(\g_reduce0[14].adder.a[14] ),
    .CO(_21308_),
    .S(_21309_));
 HA_X1 _41624_ (.A(_14074_),
    .B(_14075_),
    .CO(_21310_),
    .S(_21311_));
 HA_X1 _41625_ (.A(_14075_),
    .B(_14079_),
    .CO(_21312_),
    .S(_21313_));
 HA_X1 _41626_ (.A(_21314_),
    .B(_21315_),
    .CO(_21316_),
    .S(_21317_));
 HA_X1 _41627_ (.A(_21318_),
    .B(_21319_),
    .CO(_21320_),
    .S(_21321_));
 HA_X1 _41628_ (.A(_21322_),
    .B(_21319_),
    .CO(_21323_),
    .S(_21324_));
 HA_X1 _41629_ (.A(_21325_),
    .B(_21326_),
    .CO(_21327_),
    .S(_21328_));
 HA_X1 _41630_ (.A(_21329_),
    .B(_21326_),
    .CO(_21330_),
    .S(_21331_));
 HA_X1 _41631_ (.A(_21332_),
    .B(_21333_),
    .CO(_21334_),
    .S(_21335_));
 HA_X1 _41632_ (.A(_21336_),
    .B(_21333_),
    .CO(_21337_),
    .S(_21338_));
 HA_X1 _41633_ (.A(_21339_),
    .B(_21340_),
    .CO(_21341_),
    .S(_21342_));
 HA_X1 _41634_ (.A(_21343_),
    .B(_21340_),
    .CO(_21344_),
    .S(_21345_));
 HA_X1 _41635_ (.A(_21346_),
    .B(_21347_),
    .CO(_21348_),
    .S(_21349_));
 HA_X1 _41636_ (.A(_21350_),
    .B(_21347_),
    .CO(_21351_),
    .S(_21352_));
 HA_X1 _41637_ (.A(_21353_),
    .B(_21354_),
    .CO(_21355_),
    .S(_21356_));
 HA_X1 _41638_ (.A(_21357_),
    .B(_21354_),
    .CO(_21358_),
    .S(_21359_));
 HA_X1 _41639_ (.A(_21315_),
    .B(_21360_),
    .CO(_21361_),
    .S(_21362_));
 HA_X1 _41640_ (.A(_21363_),
    .B(_21364_),
    .CO(_21365_),
    .S(_21366_));
 HA_X1 _41641_ (.A(_21367_),
    .B(_21364_),
    .CO(_21368_),
    .S(_21369_));
 HA_X1 _41642_ (.A(_21370_),
    .B(_21371_),
    .CO(_14073_),
    .S(_21372_));
 HA_X1 _41643_ (.A(_21371_),
    .B(_21373_),
    .CO(_14078_),
    .S(_21374_));
 HA_X1 _41644_ (.A(_21375_),
    .B(_21376_),
    .CO(_21377_),
    .S(_14083_));
 HA_X1 _41645_ (.A(_21378_),
    .B(_21376_),
    .CO(_21379_),
    .S(_21380_));
 HA_X1 _41646_ (.A(_21378_),
    .B(_21376_),
    .CO(_21381_),
    .S(_21382_));
 HA_X1 _41647_ (.A(_21383_),
    .B(_21384_),
    .CO(_21385_),
    .S(_21386_));
 HA_X1 _41648_ (.A(_21375_),
    .B(_21387_),
    .CO(_14087_),
    .S(_21388_));
 HA_X1 _41649_ (.A(_21389_),
    .B(_21390_),
    .CO(_21391_),
    .S(_21392_));
 HA_X1 _41650_ (.A(_21393_),
    .B(_14082_),
    .CO(_21394_),
    .S(_21395_));
 HA_X1 _41651_ (.A(_14082_),
    .B(_14083_),
    .CO(_21396_),
    .S(_21397_));
 HA_X1 _41652_ (.A(_21398_),
    .B(_21391_),
    .CO(_21399_),
    .S(_21400_));
 HA_X1 _41653_ (.A(_21401_),
    .B(_21402_),
    .CO(_21403_),
    .S(_21404_));
 HA_X1 _41654_ (.A(_21405_),
    .B(_21406_),
    .CO(_21407_),
    .S(_21408_));
 HA_X1 _41655_ (.A(_21409_),
    .B(\g_reduce0[2].adder.a[13] ),
    .CO(_21410_),
    .S(_21411_));
 HA_X1 _41656_ (.A(_21412_),
    .B(\g_reduce0[2].adder.a[12] ),
    .CO(_21413_),
    .S(_21414_));
 HA_X1 _41657_ (.A(_21415_),
    .B(\g_reduce0[2].adder.a[11] ),
    .CO(_21416_),
    .S(_21417_));
 HA_X1 _41658_ (.A(_21418_),
    .B(\g_reduce0[2].adder.a[9] ),
    .CO(_21419_),
    .S(_21420_));
 HA_X1 _41659_ (.A(_21421_),
    .B(\g_reduce0[2].adder.a[8] ),
    .CO(_21422_),
    .S(_21423_));
 HA_X1 _41660_ (.A(_21424_),
    .B(\g_reduce0[2].adder.a[7] ),
    .CO(_21425_),
    .S(_21426_));
 HA_X1 _41661_ (.A(_21427_),
    .B(\g_reduce0[2].adder.a[6] ),
    .CO(_21428_),
    .S(_21429_));
 HA_X1 _41662_ (.A(_21430_),
    .B(\g_reduce0[2].adder.a[5] ),
    .CO(_21431_),
    .S(_21432_));
 HA_X1 _41663_ (.A(_21433_),
    .B(\g_reduce0[2].adder.a[4] ),
    .CO(_21434_),
    .S(_21435_));
 HA_X1 _41664_ (.A(_21436_),
    .B(\g_reduce0[2].adder.a[3] ),
    .CO(_21437_),
    .S(_21438_));
 HA_X1 _41665_ (.A(_21439_),
    .B(\g_reduce0[2].adder.a[2] ),
    .CO(_21440_),
    .S(_21441_));
 HA_X1 _41666_ (.A(_21442_),
    .B(\g_reduce0[2].adder.a[1] ),
    .CO(_21443_),
    .S(_21444_));
 HA_X1 _41667_ (.A(\g_reduce0[2].adder.b[0] ),
    .B(_21445_),
    .CO(_21446_),
    .S(_21447_));
 HA_X1 _41668_ (.A(\g_reduce0[2].adder.b[10] ),
    .B(_21448_),
    .CO(_21449_),
    .S(_21450_));
 HA_X1 _41669_ (.A(_21417_),
    .B(_21451_),
    .CO(_21452_),
    .S(_21453_));
 HA_X1 _41670_ (.A(_21454_),
    .B(\g_reduce0[2].adder.a[14] ),
    .CO(_21455_),
    .S(_21456_));
 HA_X1 _41671_ (.A(_14089_),
    .B(_14090_),
    .CO(_21457_),
    .S(_21458_));
 HA_X1 _41672_ (.A(_14090_),
    .B(_14094_),
    .CO(_21459_),
    .S(_21460_));
 HA_X1 _41673_ (.A(_21461_),
    .B(_21462_),
    .CO(_21463_),
    .S(_21464_));
 HA_X1 _41674_ (.A(_21465_),
    .B(_21466_),
    .CO(_21467_),
    .S(_21468_));
 HA_X1 _41675_ (.A(_21469_),
    .B(_21466_),
    .CO(_21470_),
    .S(_21471_));
 HA_X1 _41676_ (.A(_21472_),
    .B(_21473_),
    .CO(_21474_),
    .S(_21475_));
 HA_X1 _41677_ (.A(_21476_),
    .B(_21473_),
    .CO(_21477_),
    .S(_21478_));
 HA_X1 _41678_ (.A(_21479_),
    .B(_21480_),
    .CO(_21481_),
    .S(_21482_));
 HA_X1 _41679_ (.A(_21483_),
    .B(_21480_),
    .CO(_21484_),
    .S(_21485_));
 HA_X1 _41680_ (.A(_21486_),
    .B(_21487_),
    .CO(_21488_),
    .S(_21489_));
 HA_X1 _41681_ (.A(_21490_),
    .B(_21487_),
    .CO(_21491_),
    .S(_21492_));
 HA_X1 _41682_ (.A(_21493_),
    .B(_21494_),
    .CO(_21495_),
    .S(_21496_));
 HA_X1 _41683_ (.A(_21497_),
    .B(_21494_),
    .CO(_21498_),
    .S(_21499_));
 HA_X1 _41684_ (.A(_21500_),
    .B(_21501_),
    .CO(_21502_),
    .S(_21503_));
 HA_X1 _41685_ (.A(_21504_),
    .B(_21501_),
    .CO(_21505_),
    .S(_21506_));
 HA_X1 _41686_ (.A(_21462_),
    .B(_21507_),
    .CO(_21508_),
    .S(_21509_));
 HA_X1 _41687_ (.A(_21510_),
    .B(_21511_),
    .CO(_21512_),
    .S(_21513_));
 HA_X1 _41688_ (.A(_21514_),
    .B(_21511_),
    .CO(_21515_),
    .S(_21516_));
 HA_X1 _41689_ (.A(_21517_),
    .B(_21518_),
    .CO(_14088_),
    .S(_21519_));
 HA_X1 _41690_ (.A(_21518_),
    .B(_21520_),
    .CO(_14093_),
    .S(_21521_));
 HA_X1 _41691_ (.A(_21522_),
    .B(_21523_),
    .CO(_21524_),
    .S(_14098_));
 HA_X1 _41692_ (.A(_21522_),
    .B(_21525_),
    .CO(_21526_),
    .S(_21527_));
 HA_X1 _41693_ (.A(_21522_),
    .B(_21525_),
    .CO(_21528_),
    .S(_21529_));
 HA_X1 _41694_ (.A(_21530_),
    .B(_21531_),
    .CO(_21532_),
    .S(_21533_));
 HA_X1 _41695_ (.A(_21534_),
    .B(_21523_),
    .CO(_14102_),
    .S(_21535_));
 HA_X1 _41696_ (.A(_21536_),
    .B(_21537_),
    .CO(_21538_),
    .S(_21539_));
 HA_X1 _41697_ (.A(_21540_),
    .B(_14097_),
    .CO(_21541_),
    .S(_21542_));
 HA_X1 _41698_ (.A(_14097_),
    .B(_14098_),
    .CO(_21543_),
    .S(_21544_));
 HA_X1 _41699_ (.A(_21545_),
    .B(_21538_),
    .CO(_21546_),
    .S(_21547_));
 HA_X1 _41700_ (.A(_21548_),
    .B(_21549_),
    .CO(_21550_),
    .S(_21551_));
 HA_X1 _41701_ (.A(_21552_),
    .B(_21553_),
    .CO(_21554_),
    .S(_21555_));
 HA_X1 _41702_ (.A(\g_reduce0[4].adder.b[13] ),
    .B(_21556_),
    .CO(_21557_),
    .S(_21558_));
 HA_X1 _41703_ (.A(\g_reduce0[4].adder.b[12] ),
    .B(_21559_),
    .CO(_21560_),
    .S(_21561_));
 HA_X1 _41704_ (.A(\g_reduce0[4].adder.b[11] ),
    .B(_21562_),
    .CO(_21563_),
    .S(_21564_));
 HA_X1 _41705_ (.A(_21565_),
    .B(\g_reduce0[4].adder.a[10] ),
    .CO(_21566_),
    .S(_21567_));
 HA_X1 _41706_ (.A(\g_reduce0[4].adder.b[9] ),
    .B(_21568_),
    .CO(_21569_),
    .S(_21570_));
 HA_X1 _41707_ (.A(\g_reduce0[4].adder.b[8] ),
    .B(_21571_),
    .CO(_21572_),
    .S(_21573_));
 HA_X1 _41708_ (.A(\g_reduce0[4].adder.b[7] ),
    .B(_21574_),
    .CO(_21575_),
    .S(_21576_));
 HA_X1 _41709_ (.A(\g_reduce0[4].adder.b[6] ),
    .B(_21577_),
    .CO(_21578_),
    .S(_21579_));
 HA_X1 _41710_ (.A(\g_reduce0[4].adder.b[5] ),
    .B(_21580_),
    .CO(_21581_),
    .S(_21582_));
 HA_X1 _41711_ (.A(\g_reduce0[4].adder.b[4] ),
    .B(_21583_),
    .CO(_21584_),
    .S(_21585_));
 HA_X1 _41712_ (.A(\g_reduce0[4].adder.b[3] ),
    .B(_21586_),
    .CO(_21587_),
    .S(_21588_));
 HA_X1 _41713_ (.A(\g_reduce0[4].adder.b[2] ),
    .B(_21589_),
    .CO(_21590_),
    .S(_21591_));
 HA_X1 _41714_ (.A(\g_reduce0[4].adder.b[1] ),
    .B(_21592_),
    .CO(_21593_),
    .S(_21594_));
 HA_X1 _41715_ (.A(_21595_),
    .B(_21564_),
    .CO(_21596_),
    .S(_21597_));
 HA_X1 _41716_ (.A(\g_reduce0[4].adder.b[14] ),
    .B(_21598_),
    .CO(_21599_),
    .S(_21600_));
 HA_X1 _41717_ (.A(_14104_),
    .B(_14105_),
    .CO(_21601_),
    .S(_21602_));
 HA_X1 _41718_ (.A(_14105_),
    .B(_14109_),
    .CO(_21603_),
    .S(_21604_));
 HA_X1 _41719_ (.A(_21605_),
    .B(_21606_),
    .CO(_21607_),
    .S(_21608_));
 HA_X1 _41720_ (.A(_21609_),
    .B(_21610_),
    .CO(_21611_),
    .S(_21612_));
 HA_X1 _41721_ (.A(_21613_),
    .B(_21610_),
    .CO(_21614_),
    .S(_21615_));
 HA_X1 _41722_ (.A(_21616_),
    .B(_21617_),
    .CO(_21618_),
    .S(_21619_));
 HA_X1 _41723_ (.A(_21620_),
    .B(_21617_),
    .CO(_21621_),
    .S(_21622_));
 HA_X1 _41724_ (.A(_21623_),
    .B(_21624_),
    .CO(_21625_),
    .S(_21626_));
 HA_X1 _41725_ (.A(_21627_),
    .B(_21624_),
    .CO(_21628_),
    .S(_21629_));
 HA_X1 _41726_ (.A(_21630_),
    .B(_21631_),
    .CO(_21632_),
    .S(_21633_));
 HA_X1 _41727_ (.A(_21634_),
    .B(_21631_),
    .CO(_21635_),
    .S(_21636_));
 HA_X1 _41728_ (.A(_21637_),
    .B(_21638_),
    .CO(_21639_),
    .S(_21640_));
 HA_X1 _41729_ (.A(_21641_),
    .B(_21638_),
    .CO(_21642_),
    .S(_21643_));
 HA_X1 _41730_ (.A(_21644_),
    .B(_21645_),
    .CO(_21646_),
    .S(_21647_));
 HA_X1 _41731_ (.A(_21648_),
    .B(_21645_),
    .CO(_21649_),
    .S(_21650_));
 HA_X1 _41732_ (.A(_21651_),
    .B(_21606_),
    .CO(_21652_),
    .S(_21653_));
 HA_X1 _41733_ (.A(_21654_),
    .B(_21655_),
    .CO(_21656_),
    .S(_21657_));
 HA_X1 _41734_ (.A(_21654_),
    .B(_21658_),
    .CO(_21659_),
    .S(_21660_));
 HA_X1 _41735_ (.A(_21661_),
    .B(_21662_),
    .CO(_14103_),
    .S(_21663_));
 HA_X1 _41736_ (.A(_21662_),
    .B(_21664_),
    .CO(_14108_),
    .S(_21665_));
 HA_X1 _41737_ (.A(_21666_),
    .B(_21667_),
    .CO(_21668_),
    .S(_14112_));
 HA_X1 _41738_ (.A(_21669_),
    .B(_21667_),
    .CO(_21670_),
    .S(_21671_));
 HA_X1 _41739_ (.A(_21669_),
    .B(_21667_),
    .CO(_21672_),
    .S(_21673_));
 HA_X1 _41740_ (.A(_21674_),
    .B(_21675_),
    .CO(_21676_),
    .S(_21677_));
 HA_X1 _41741_ (.A(_21666_),
    .B(_21678_),
    .CO(_14117_),
    .S(_21679_));
 HA_X1 _41742_ (.A(_21680_),
    .B(_21681_),
    .CO(_21682_),
    .S(_21683_));
 HA_X1 _41743_ (.A(_21684_),
    .B(_14113_),
    .CO(_21685_),
    .S(_21686_));
 HA_X1 _41744_ (.A(_14112_),
    .B(_14113_),
    .CO(_21687_),
    .S(_21688_));
 HA_X1 _41745_ (.A(_21689_),
    .B(_21682_),
    .CO(_21690_),
    .S(_21691_));
 HA_X1 _41746_ (.A(_21692_),
    .B(_21693_),
    .CO(_21694_),
    .S(_21695_));
 HA_X1 _41747_ (.A(_21696_),
    .B(_21697_),
    .CO(_21698_),
    .S(_21699_));
 HA_X1 _41748_ (.A(_21700_),
    .B(\g_reduce0[6].adder.a[13] ),
    .CO(_21701_),
    .S(_21702_));
 HA_X1 _41749_ (.A(_21703_),
    .B(\g_reduce0[6].adder.a[12] ),
    .CO(_21704_),
    .S(_21705_));
 HA_X1 _41750_ (.A(_21706_),
    .B(\g_reduce0[6].adder.a[11] ),
    .CO(_21707_),
    .S(_21708_));
 HA_X1 _41751_ (.A(_21709_),
    .B(\g_reduce0[6].adder.a[9] ),
    .CO(_21710_),
    .S(_21711_));
 HA_X1 _41752_ (.A(_21712_),
    .B(\g_reduce0[6].adder.a[8] ),
    .CO(_21713_),
    .S(_21714_));
 HA_X1 _41753_ (.A(_21715_),
    .B(\g_reduce0[6].adder.a[7] ),
    .CO(_21716_),
    .S(_21717_));
 HA_X1 _41754_ (.A(_21718_),
    .B(\g_reduce0[6].adder.a[6] ),
    .CO(_21719_),
    .S(_21720_));
 HA_X1 _41755_ (.A(_21721_),
    .B(\g_reduce0[6].adder.a[5] ),
    .CO(_21722_),
    .S(_21723_));
 HA_X1 _41756_ (.A(_21724_),
    .B(\g_reduce0[6].adder.a[4] ),
    .CO(_21725_),
    .S(_21726_));
 HA_X1 _41757_ (.A(_21727_),
    .B(\g_reduce0[6].adder.a[3] ),
    .CO(_21728_),
    .S(_21729_));
 HA_X1 _41758_ (.A(_21730_),
    .B(\g_reduce0[6].adder.a[2] ),
    .CO(_21731_),
    .S(_21732_));
 HA_X1 _41759_ (.A(_21733_),
    .B(\g_reduce0[6].adder.a[1] ),
    .CO(_21734_),
    .S(_21735_));
 HA_X1 _41760_ (.A(\g_reduce0[6].adder.b[0] ),
    .B(_21736_),
    .CO(_21737_),
    .S(_21738_));
 HA_X1 _41761_ (.A(\g_reduce0[6].adder.b[10] ),
    .B(_21739_),
    .CO(_21740_),
    .S(_21741_));
 HA_X1 _41762_ (.A(_21742_),
    .B(_21708_),
    .CO(_21743_),
    .S(_21744_));
 HA_X1 _41763_ (.A(_21745_),
    .B(\g_reduce0[6].adder.a[14] ),
    .CO(_21746_),
    .S(_21747_));
 HA_X1 _41764_ (.A(_14119_),
    .B(_14120_),
    .CO(_21748_),
    .S(_21749_));
 HA_X1 _41765_ (.A(_14120_),
    .B(_14124_),
    .CO(_21750_),
    .S(_21751_));
 HA_X1 _41766_ (.A(_21752_),
    .B(_21753_),
    .CO(_21754_),
    .S(_21755_));
 HA_X1 _41767_ (.A(_21756_),
    .B(_21757_),
    .CO(_21758_),
    .S(_21759_));
 HA_X1 _41768_ (.A(_21760_),
    .B(_21757_),
    .CO(_21761_),
    .S(_21762_));
 HA_X1 _41769_ (.A(_21763_),
    .B(_21764_),
    .CO(_21765_),
    .S(_21766_));
 HA_X1 _41770_ (.A(_21767_),
    .B(_21764_),
    .CO(_21768_),
    .S(_21769_));
 HA_X1 _41771_ (.A(_21770_),
    .B(_21771_),
    .CO(_21772_),
    .S(_21773_));
 HA_X1 _41772_ (.A(_21774_),
    .B(_21771_),
    .CO(_21775_),
    .S(_21776_));
 HA_X1 _41773_ (.A(_21777_),
    .B(_21778_),
    .CO(_21779_),
    .S(_21780_));
 HA_X1 _41774_ (.A(_21781_),
    .B(_21778_),
    .CO(_21782_),
    .S(_21783_));
 HA_X1 _41775_ (.A(_21784_),
    .B(_21785_),
    .CO(_21786_),
    .S(_21787_));
 HA_X1 _41776_ (.A(_21788_),
    .B(_21785_),
    .CO(_21789_),
    .S(_21790_));
 HA_X1 _41777_ (.A(_21791_),
    .B(_21792_),
    .CO(_21793_),
    .S(_21794_));
 HA_X1 _41778_ (.A(_21795_),
    .B(_21792_),
    .CO(_21796_),
    .S(_21797_));
 HA_X1 _41779_ (.A(_21753_),
    .B(_21798_),
    .CO(_21799_),
    .S(_21800_));
 HA_X1 _41780_ (.A(_21801_),
    .B(_21802_),
    .CO(_21803_),
    .S(_21804_));
 HA_X1 _41781_ (.A(_21805_),
    .B(_21802_),
    .CO(_21806_),
    .S(_21807_));
 HA_X1 _41782_ (.A(_21808_),
    .B(_21809_),
    .CO(_14118_),
    .S(_21810_));
 HA_X1 _41783_ (.A(_21809_),
    .B(_21811_),
    .CO(_14123_),
    .S(_21812_));
 HA_X1 _41784_ (.A(_21813_),
    .B(_21814_),
    .CO(_21815_),
    .S(_14128_));
 HA_X1 _41785_ (.A(_21813_),
    .B(_21816_),
    .CO(_21817_),
    .S(_21818_));
 HA_X1 _41786_ (.A(_21813_),
    .B(_21816_),
    .CO(_21819_),
    .S(_21820_));
 HA_X1 _41787_ (.A(_21821_),
    .B(_21822_),
    .CO(_21823_),
    .S(_21824_));
 HA_X1 _41788_ (.A(_21825_),
    .B(_21814_),
    .CO(_14132_),
    .S(_21826_));
 HA_X1 _41789_ (.A(_21827_),
    .B(_21828_),
    .CO(_21829_),
    .S(_21830_));
 HA_X1 _41790_ (.A(_21831_),
    .B(_14127_),
    .CO(_21832_),
    .S(_21833_));
 HA_X1 _41791_ (.A(_14127_),
    .B(_14128_),
    .CO(_21834_),
    .S(_21835_));
 HA_X1 _41792_ (.A(_21836_),
    .B(_21829_),
    .CO(_21837_),
    .S(_21838_));
 HA_X1 _41793_ (.A(_21839_),
    .B(_21840_),
    .CO(_21841_),
    .S(_21842_));
 HA_X1 _41794_ (.A(_21843_),
    .B(_21844_),
    .CO(_21845_),
    .S(_21846_));
 HA_X1 _41795_ (.A(\g_reduce0[8].adder.b[13] ),
    .B(_21847_),
    .CO(_21848_),
    .S(_21849_));
 HA_X1 _41796_ (.A(\g_reduce0[8].adder.b[12] ),
    .B(_21850_),
    .CO(_21851_),
    .S(_21852_));
 HA_X1 _41797_ (.A(\g_reduce0[8].adder.b[11] ),
    .B(_21853_),
    .CO(_21854_),
    .S(_21855_));
 HA_X1 _41798_ (.A(_21856_),
    .B(\g_reduce0[8].adder.a[10] ),
    .CO(_21857_),
    .S(_21858_));
 HA_X1 _41799_ (.A(\g_reduce0[8].adder.b[9] ),
    .B(_21859_),
    .CO(_21860_),
    .S(_21861_));
 HA_X1 _41800_ (.A(\g_reduce0[8].adder.b[8] ),
    .B(_21862_),
    .CO(_21863_),
    .S(_21864_));
 HA_X1 _41801_ (.A(\g_reduce0[8].adder.b[7] ),
    .B(_21865_),
    .CO(_21866_),
    .S(_21867_));
 HA_X1 _41802_ (.A(\g_reduce0[8].adder.b[6] ),
    .B(_21868_),
    .CO(_21869_),
    .S(_21870_));
 HA_X1 _41803_ (.A(\g_reduce0[8].adder.b[5] ),
    .B(_21871_),
    .CO(_21872_),
    .S(_21873_));
 HA_X1 _41804_ (.A(\g_reduce0[8].adder.b[4] ),
    .B(_21874_),
    .CO(_21875_),
    .S(_21876_));
 HA_X1 _41805_ (.A(\g_reduce0[8].adder.b[3] ),
    .B(_21877_),
    .CO(_21878_),
    .S(_21879_));
 HA_X1 _41806_ (.A(\g_reduce0[8].adder.b[2] ),
    .B(_21880_),
    .CO(_21881_),
    .S(_21882_));
 HA_X1 _41807_ (.A(\g_reduce0[8].adder.b[1] ),
    .B(_21883_),
    .CO(_21884_),
    .S(_21885_));
 HA_X1 _41808_ (.A(_21855_),
    .B(_21886_),
    .CO(_21887_),
    .S(_21888_));
 HA_X1 _41809_ (.A(\g_reduce0[8].adder.b[14] ),
    .B(_21889_),
    .CO(_21890_),
    .S(_21891_));
 HA_X1 _41810_ (.A(_14133_),
    .B(_14134_),
    .CO(_21892_),
    .S(_21893_));
 HA_X1 _41811_ (.A(_14134_),
    .B(_14139_),
    .CO(_21894_),
    .S(_21895_));
 HA_X1 _41812_ (.A(_21896_),
    .B(_21897_),
    .CO(_21898_),
    .S(_21899_));
 HA_X1 _41813_ (.A(_21900_),
    .B(_21901_),
    .CO(_21902_),
    .S(_21903_));
 HA_X1 _41814_ (.A(_21904_),
    .B(_21901_),
    .CO(_21905_),
    .S(_21906_));
 HA_X1 _41815_ (.A(_21907_),
    .B(_21908_),
    .CO(_21909_),
    .S(_21910_));
 HA_X1 _41816_ (.A(_21911_),
    .B(_21908_),
    .CO(_21912_),
    .S(_21913_));
 HA_X1 _41817_ (.A(_21914_),
    .B(_21915_),
    .CO(_21916_),
    .S(_21917_));
 HA_X1 _41818_ (.A(_21918_),
    .B(_21915_),
    .CO(_21919_),
    .S(_21920_));
 HA_X1 _41819_ (.A(_21921_),
    .B(_21922_),
    .CO(_21923_),
    .S(_21924_));
 HA_X1 _41820_ (.A(_21925_),
    .B(_21922_),
    .CO(_21926_),
    .S(_21927_));
 HA_X1 _41821_ (.A(_21928_),
    .B(_21929_),
    .CO(_21930_),
    .S(_21931_));
 HA_X1 _41822_ (.A(_21932_),
    .B(_21929_),
    .CO(_21933_),
    .S(_21934_));
 HA_X1 _41823_ (.A(_21935_),
    .B(_21936_),
    .CO(_21937_),
    .S(_21938_));
 HA_X1 _41824_ (.A(_21939_),
    .B(_21936_),
    .CO(_21940_),
    .S(_21941_));
 HA_X1 _41825_ (.A(_21942_),
    .B(_21897_),
    .CO(_21943_),
    .S(_21944_));
 HA_X1 _41826_ (.A(_21945_),
    .B(_21946_),
    .CO(_21947_),
    .S(_21948_));
 HA_X1 _41827_ (.A(_21949_),
    .B(_21946_),
    .CO(_21950_),
    .S(_21951_));
 HA_X1 _41828_ (.A(_21952_),
    .B(_21953_),
    .CO(_14135_),
    .S(_21954_));
 HA_X1 _41829_ (.A(_21955_),
    .B(_21953_),
    .CO(_14138_),
    .S(_21956_));
 HA_X1 _41830_ (.A(_21957_),
    .B(_21958_),
    .CO(_21959_),
    .S(_14143_));
 HA_X1 _41831_ (.A(_21957_),
    .B(_21960_),
    .CO(_21961_),
    .S(_21962_));
 HA_X1 _41832_ (.A(_21957_),
    .B(_21960_),
    .CO(_21963_),
    .S(_21964_));
 HA_X1 _41833_ (.A(_21965_),
    .B(_21966_),
    .CO(_21967_),
    .S(_21968_));
 HA_X1 _41834_ (.A(_21958_),
    .B(_21969_),
    .CO(_14147_),
    .S(_21970_));
 HA_X1 _41835_ (.A(_21971_),
    .B(_21972_),
    .CO(_21973_),
    .S(_21974_));
 HA_X1 _41836_ (.A(_21975_),
    .B(_14144_),
    .CO(_21976_),
    .S(_21977_));
 HA_X1 _41837_ (.A(_14143_),
    .B(_14144_),
    .CO(_21978_),
    .S(_21979_));
 HA_X1 _41838_ (.A(_21980_),
    .B(_21973_),
    .CO(_21981_),
    .S(_21982_));
 HA_X1 _41839_ (.A(_21983_),
    .B(_21984_),
    .CO(_21985_),
    .S(_21986_));
 HA_X1 _41840_ (.A(_21987_),
    .B(_21988_),
    .CO(_21989_),
    .S(_21990_));
 HA_X1 _41841_ (.A(_21991_),
    .B(\g_reduce0[2].adder.x[13] ),
    .CO(_21992_),
    .S(_21993_));
 HA_X1 _41842_ (.A(_21994_),
    .B(\g_reduce0[2].adder.x[12] ),
    .CO(_21995_),
    .S(_21996_));
 HA_X1 _41843_ (.A(_21997_),
    .B(\g_reduce0[2].adder.x[11] ),
    .CO(_21998_),
    .S(_21999_));
 HA_X1 _41844_ (.A(\g_reduce0[0].adder.x[10] ),
    .B(_22000_),
    .CO(_22001_),
    .S(_22002_));
 HA_X1 _41845_ (.A(_22003_),
    .B(\g_reduce0[2].adder.x[9] ),
    .CO(_22004_),
    .S(_22005_));
 HA_X1 _41846_ (.A(_22006_),
    .B(\g_reduce0[2].adder.x[8] ),
    .CO(_22007_),
    .S(_22008_));
 HA_X1 _41847_ (.A(_22009_),
    .B(\g_reduce0[2].adder.x[7] ),
    .CO(_22010_),
    .S(_22011_));
 HA_X1 _41848_ (.A(_22012_),
    .B(\g_reduce0[2].adder.x[6] ),
    .CO(_22013_),
    .S(_22014_));
 HA_X1 _41849_ (.A(_22015_),
    .B(\g_reduce0[2].adder.x[5] ),
    .CO(_22016_),
    .S(_22017_));
 HA_X1 _41850_ (.A(_22018_),
    .B(\g_reduce0[2].adder.x[4] ),
    .CO(_22019_),
    .S(_22020_));
 HA_X1 _41851_ (.A(_22021_),
    .B(\g_reduce0[2].adder.x[3] ),
    .CO(_22022_),
    .S(_22023_));
 HA_X1 _41852_ (.A(_22024_),
    .B(\g_reduce0[2].adder.x[2] ),
    .CO(_22025_),
    .S(_22026_));
 HA_X1 _41853_ (.A(_22027_),
    .B(\g_reduce0[2].adder.x[1] ),
    .CO(_22028_),
    .S(_22029_));
 HA_X1 _41854_ (.A(_21999_),
    .B(_22030_),
    .CO(_22031_),
    .S(_22032_));
 HA_X1 _41855_ (.A(_22033_),
    .B(\g_reduce0[2].adder.x[14] ),
    .CO(_22034_),
    .S(_22035_));
 HA_X1 _41856_ (.A(_14148_),
    .B(_14149_),
    .CO(_22036_),
    .S(_22037_));
 HA_X1 _41857_ (.A(_14148_),
    .B(_14153_),
    .CO(_22038_),
    .S(_22039_));
 HA_X1 _41858_ (.A(_22040_),
    .B(_22041_),
    .CO(_22042_),
    .S(_22043_));
 HA_X1 _41859_ (.A(_22044_),
    .B(_22045_),
    .CO(_22046_),
    .S(_22047_));
 HA_X1 _41860_ (.A(_22044_),
    .B(_22048_),
    .CO(_22049_),
    .S(_22050_));
 HA_X1 _41861_ (.A(_22051_),
    .B(_22052_),
    .CO(_22053_),
    .S(_22054_));
 HA_X1 _41862_ (.A(_22051_),
    .B(_22055_),
    .CO(_22056_),
    .S(_22057_));
 HA_X1 _41863_ (.A(_22058_),
    .B(_22059_),
    .CO(_22060_),
    .S(_22061_));
 HA_X1 _41864_ (.A(_22058_),
    .B(_22062_),
    .CO(_22063_),
    .S(_22064_));
 HA_X1 _41865_ (.A(_22065_),
    .B(_22066_),
    .CO(_22067_),
    .S(_22068_));
 HA_X1 _41866_ (.A(_22065_),
    .B(_22069_),
    .CO(_22070_),
    .S(_22071_));
 HA_X1 _41867_ (.A(_22072_),
    .B(_22073_),
    .CO(_22074_),
    .S(_22075_));
 HA_X1 _41868_ (.A(_22072_),
    .B(_22076_),
    .CO(_22077_),
    .S(_22078_));
 HA_X1 _41869_ (.A(_22079_),
    .B(_22080_),
    .CO(_22081_),
    .S(_22082_));
 HA_X1 _41870_ (.A(_22083_),
    .B(_22080_),
    .CO(_22084_),
    .S(_22085_));
 HA_X1 _41871_ (.A(_22086_),
    .B(_22041_),
    .CO(_22087_),
    .S(_22088_));
 HA_X1 _41872_ (.A(_22089_),
    .B(_22090_),
    .CO(_22091_),
    .S(_22092_));
 HA_X1 _41873_ (.A(_22089_),
    .B(_22093_),
    .CO(_22094_),
    .S(_22095_));
 HA_X1 _41874_ (.A(_22096_),
    .B(_22097_),
    .CO(_14150_),
    .S(_22098_));
 HA_X1 _41875_ (.A(_22099_),
    .B(_22097_),
    .CO(_14154_),
    .S(_22100_));
 HA_X1 _41876_ (.A(_22101_),
    .B(_22102_),
    .CO(_22103_),
    .S(_14162_));
 HA_X1 _41877_ (.A(_22104_),
    .B(_22102_),
    .CO(_22105_),
    .S(_22106_));
 HA_X1 _41878_ (.A(_22104_),
    .B(_22102_),
    .CO(_22107_),
    .S(_22108_));
 HA_X1 _41879_ (.A(_22109_),
    .B(_22110_),
    .CO(_22111_),
    .S(_22112_));
 HA_X1 _41880_ (.A(_22101_),
    .B(_22113_),
    .CO(_14158_),
    .S(_22114_));
 HA_X1 _41881_ (.A(_22115_),
    .B(_22116_),
    .CO(_22117_),
    .S(_22118_));
 HA_X1 _41882_ (.A(_22119_),
    .B(_14163_),
    .CO(_22120_),
    .S(_22121_));
 HA_X1 _41883_ (.A(_14162_),
    .B(_14163_),
    .CO(_22122_),
    .S(_22123_));
 HA_X1 _41884_ (.A(_22124_),
    .B(_22117_),
    .CO(_22125_),
    .S(_22126_));
 HA_X1 _41885_ (.A(_22127_),
    .B(_22128_),
    .CO(_22129_),
    .S(_22130_));
 HA_X1 _41886_ (.A(_22131_),
    .B(_22132_),
    .CO(_22133_),
    .S(_22134_));
 HA_X1 _41887_ (.A(\g_reduce0[4].adder.x[13] ),
    .B(_22135_),
    .CO(_22136_),
    .S(_22137_));
 HA_X1 _41888_ (.A(\g_reduce0[4].adder.x[12] ),
    .B(_22138_),
    .CO(_22139_),
    .S(_22140_));
 HA_X1 _41889_ (.A(\g_reduce0[4].adder.x[11] ),
    .B(_22141_),
    .CO(_22142_),
    .S(_22143_));
 HA_X1 _41890_ (.A(\g_reduce0[4].adder.x[9] ),
    .B(_22144_),
    .CO(_22145_),
    .S(_22146_));
 HA_X1 _41891_ (.A(\g_reduce0[4].adder.x[8] ),
    .B(_22147_),
    .CO(_22148_),
    .S(_22149_));
 HA_X1 _41892_ (.A(\g_reduce0[4].adder.x[7] ),
    .B(_22150_),
    .CO(_22151_),
    .S(_22152_));
 HA_X1 _41893_ (.A(\g_reduce0[4].adder.x[6] ),
    .B(_22153_),
    .CO(_22154_),
    .S(_22155_));
 HA_X1 _41894_ (.A(\g_reduce0[4].adder.x[5] ),
    .B(_22156_),
    .CO(_22157_),
    .S(_22158_));
 HA_X1 _41895_ (.A(\g_reduce0[4].adder.x[4] ),
    .B(_22159_),
    .CO(_22160_),
    .S(_22161_));
 HA_X1 _41896_ (.A(\g_reduce0[4].adder.x[3] ),
    .B(_22162_),
    .CO(_22163_),
    .S(_22164_));
 HA_X1 _41897_ (.A(\g_reduce0[4].adder.x[2] ),
    .B(_22165_),
    .CO(_22166_),
    .S(_22167_));
 HA_X1 _41898_ (.A(\g_reduce0[4].adder.x[1] ),
    .B(_22168_),
    .CO(_22169_),
    .S(_22170_));
 HA_X1 _41899_ (.A(_22171_),
    .B(\g_reduce0[6].adder.x[0] ),
    .CO(_22172_),
    .S(_22173_));
 HA_X1 _41900_ (.A(_22174_),
    .B(\g_reduce0[6].adder.x[10] ),
    .CO(_22175_),
    .S(_22176_));
 HA_X1 _41901_ (.A(_22143_),
    .B(_22177_),
    .CO(_22178_),
    .S(_22179_));
 HA_X1 _41902_ (.A(\g_reduce0[4].adder.x[14] ),
    .B(_22180_),
    .CO(_22181_),
    .S(_22182_));
 HA_X1 _41903_ (.A(_14164_),
    .B(_14165_),
    .CO(_22183_),
    .S(_22184_));
 HA_X1 _41904_ (.A(_14165_),
    .B(_14169_),
    .CO(_22185_),
    .S(_22186_));
 HA_X1 _41905_ (.A(_22187_),
    .B(_22188_),
    .CO(_22189_),
    .S(_22190_));
 HA_X1 _41906_ (.A(_22191_),
    .B(_22192_),
    .CO(_22193_),
    .S(_22194_));
 HA_X1 _41907_ (.A(_22191_),
    .B(_22195_),
    .CO(_22196_),
    .S(_22197_));
 HA_X1 _41908_ (.A(_22198_),
    .B(_22199_),
    .CO(_22200_),
    .S(_22201_));
 HA_X1 _41909_ (.A(_22202_),
    .B(_22199_),
    .CO(_22203_),
    .S(_22204_));
 HA_X1 _41910_ (.A(_22205_),
    .B(_22206_),
    .CO(_22207_),
    .S(_22208_));
 HA_X1 _41911_ (.A(_22205_),
    .B(_22209_),
    .CO(_22210_),
    .S(_22211_));
 HA_X1 _41912_ (.A(_22212_),
    .B(_22213_),
    .CO(_22214_),
    .S(_22215_));
 HA_X1 _41913_ (.A(_22212_),
    .B(_22216_),
    .CO(_22217_),
    .S(_22218_));
 HA_X1 _41914_ (.A(_22219_),
    .B(_22220_),
    .CO(_22221_),
    .S(_22222_));
 HA_X1 _41915_ (.A(_22223_),
    .B(_22220_),
    .CO(_22224_),
    .S(_22225_));
 HA_X1 _41916_ (.A(_22226_),
    .B(_22227_),
    .CO(_22228_),
    .S(_22229_));
 HA_X1 _41917_ (.A(_22230_),
    .B(_22227_),
    .CO(_22231_),
    .S(_22232_));
 HA_X1 _41918_ (.A(_22188_),
    .B(_22233_),
    .CO(_22234_),
    .S(_22235_));
 HA_X1 _41919_ (.A(_22236_),
    .B(_22237_),
    .CO(_22238_),
    .S(_22239_));
 HA_X1 _41920_ (.A(_22236_),
    .B(_22240_),
    .CO(_22241_),
    .S(_22242_));
 HA_X1 _41921_ (.A(_22243_),
    .B(_22244_),
    .CO(_14166_),
    .S(_22245_));
 HA_X1 _41922_ (.A(_22244_),
    .B(_22246_),
    .CO(_14170_),
    .S(_22247_));
 HA_X1 _41923_ (.A(_22248_),
    .B(_22249_),
    .CO(_22250_),
    .S(_14179_));
 HA_X1 _41924_ (.A(_22248_),
    .B(_22251_),
    .CO(_22252_),
    .S(_22253_));
 HA_X1 _41925_ (.A(_22248_),
    .B(_22251_),
    .CO(_22254_),
    .S(_22255_));
 HA_X1 _41926_ (.A(_22256_),
    .B(_22257_),
    .CO(_22258_),
    .S(_22259_));
 HA_X1 _41927_ (.A(_22260_),
    .B(_22249_),
    .CO(_14175_),
    .S(_22261_));
 HA_X1 _41928_ (.A(_22262_),
    .B(_22263_),
    .CO(_22264_),
    .S(_22265_));
 HA_X1 _41929_ (.A(_14178_),
    .B(_22266_),
    .CO(_22267_),
    .S(_22268_));
 HA_X1 _41930_ (.A(_14178_),
    .B(_14179_),
    .CO(_22269_),
    .S(_22270_));
 HA_X1 _41931_ (.A(_22271_),
    .B(_22264_),
    .CO(_22272_),
    .S(_22273_));
 HA_X1 _41932_ (.A(_22274_),
    .B(_22275_),
    .CO(_22276_),
    .S(_22277_));
 HA_X1 _41933_ (.A(_22278_),
    .B(_22279_),
    .CO(_22280_),
    .S(_22281_));
 HA_X1 _41934_ (.A(_22282_),
    .B(\g_reduce0[8].adder.x[13] ),
    .CO(_22283_),
    .S(_22284_));
 HA_X1 _41935_ (.A(_22285_),
    .B(\g_reduce0[8].adder.x[12] ),
    .CO(_22286_),
    .S(_22287_));
 HA_X1 _41936_ (.A(_22288_),
    .B(\g_reduce0[8].adder.x[11] ),
    .CO(_22289_),
    .S(_22290_));
 HA_X1 _41937_ (.A(_22291_),
    .B(\g_reduce0[8].adder.x[9] ),
    .CO(_22292_),
    .S(_22293_));
 HA_X1 _41938_ (.A(_22294_),
    .B(\g_reduce0[8].adder.x[8] ),
    .CO(_22295_),
    .S(_22296_));
 HA_X1 _41939_ (.A(_22297_),
    .B(\g_reduce0[8].adder.x[7] ),
    .CO(_22298_),
    .S(_22299_));
 HA_X1 _41940_ (.A(_22300_),
    .B(\g_reduce0[8].adder.x[6] ),
    .CO(_22301_),
    .S(_22302_));
 HA_X1 _41941_ (.A(_22303_),
    .B(\g_reduce0[8].adder.x[5] ),
    .CO(_22304_),
    .S(_22305_));
 HA_X1 _41942_ (.A(_22306_),
    .B(\g_reduce0[8].adder.x[4] ),
    .CO(_22307_),
    .S(_22308_));
 HA_X1 _41943_ (.A(_22309_),
    .B(\g_reduce0[8].adder.x[3] ),
    .CO(_22310_),
    .S(_22311_));
 HA_X1 _41944_ (.A(_22312_),
    .B(\g_reduce0[8].adder.x[2] ),
    .CO(_22313_),
    .S(_22314_));
 HA_X1 _41945_ (.A(_22315_),
    .B(\g_reduce0[8].adder.x[1] ),
    .CO(_22316_),
    .S(_22317_));
 HA_X1 _41946_ (.A(\g_reduce0[10].adder.x[0] ),
    .B(_22318_),
    .CO(_22319_),
    .S(_22320_));
 HA_X1 _41947_ (.A(\g_reduce0[10].adder.x[10] ),
    .B(_22321_),
    .CO(_22322_),
    .S(_22323_));
 HA_X1 _41948_ (.A(_22290_),
    .B(_22324_),
    .CO(_22325_),
    .S(_22326_));
 HA_X1 _41949_ (.A(_22327_),
    .B(\g_reduce0[8].adder.x[14] ),
    .CO(_22328_),
    .S(_22329_));
 HA_X1 _41950_ (.A(_14180_),
    .B(_14182_),
    .CO(_22330_),
    .S(_22331_));
 HA_X1 _41951_ (.A(_14182_),
    .B(_14186_),
    .CO(_22332_),
    .S(_22333_));
 HA_X1 _41952_ (.A(_22334_),
    .B(_22335_),
    .CO(_22336_),
    .S(_22337_));
 HA_X1 _41953_ (.A(_22338_),
    .B(_22339_),
    .CO(_22340_),
    .S(_22341_));
 HA_X1 _41954_ (.A(_22338_),
    .B(_22342_),
    .CO(_22343_),
    .S(_22344_));
 HA_X1 _41955_ (.A(_22345_),
    .B(_22346_),
    .CO(_22347_),
    .S(_22348_));
 HA_X1 _41956_ (.A(_22349_),
    .B(_22346_),
    .CO(_22350_),
    .S(_22351_));
 HA_X1 _41957_ (.A(_22352_),
    .B(_22353_),
    .CO(_22354_),
    .S(_22355_));
 HA_X1 _41958_ (.A(_22352_),
    .B(_22356_),
    .CO(_22357_),
    .S(_22358_));
 HA_X1 _41959_ (.A(_22359_),
    .B(_22360_),
    .CO(_22361_),
    .S(_22362_));
 HA_X1 _41960_ (.A(_22359_),
    .B(_22363_),
    .CO(_22364_),
    .S(_22365_));
 HA_X1 _41961_ (.A(_22366_),
    .B(_22367_),
    .CO(_22368_),
    .S(_22369_));
 HA_X1 _41962_ (.A(_22370_),
    .B(_22367_),
    .CO(_22371_),
    .S(_22372_));
 HA_X1 _41963_ (.A(_22373_),
    .B(_22374_),
    .CO(_22375_),
    .S(_22376_));
 HA_X1 _41964_ (.A(_22377_),
    .B(_22374_),
    .CO(_22378_),
    .S(_22379_));
 HA_X1 _41965_ (.A(_22335_),
    .B(_22380_),
    .CO(_22381_),
    .S(_22382_));
 HA_X1 _41966_ (.A(_22383_),
    .B(_22384_),
    .CO(_22385_),
    .S(_22386_));
 HA_X1 _41967_ (.A(_22387_),
    .B(_22384_),
    .CO(_22388_),
    .S(_22389_));
 HA_X1 _41968_ (.A(_22390_),
    .B(_22391_),
    .CO(_14181_),
    .S(_22392_));
 HA_X1 _41969_ (.A(_22393_),
    .B(_22391_),
    .CO(_14185_),
    .S(_22394_));
 HA_X1 _41970_ (.A(_22395_),
    .B(_22396_),
    .CO(_22397_),
    .S(_14190_));
 HA_X1 _41971_ (.A(_22395_),
    .B(_22398_),
    .CO(_22399_),
    .S(_22400_));
 HA_X1 _41972_ (.A(_22395_),
    .B(_22398_),
    .CO(_22401_),
    .S(_22402_));
 HA_X1 _41973_ (.A(_22403_),
    .B(_22404_),
    .CO(_22405_),
    .S(_22406_));
 HA_X1 _41974_ (.A(_22407_),
    .B(_22396_),
    .CO(_14194_),
    .S(_22408_));
 HA_X1 _41975_ (.A(_22409_),
    .B(_22410_),
    .CO(_22411_),
    .S(_22412_));
 HA_X1 _41976_ (.A(_22413_),
    .B(_14189_),
    .CO(_22414_),
    .S(_22415_));
 HA_X1 _41977_ (.A(_14189_),
    .B(_14190_),
    .CO(_22416_),
    .S(_22417_));
 HA_X1 _41978_ (.A(_22418_),
    .B(_22411_),
    .CO(_22419_),
    .S(_22420_));
 HA_X1 _41979_ (.A(_22421_),
    .B(_22422_),
    .CO(_22423_),
    .S(_22424_));
 HA_X1 _41980_ (.A(_22425_),
    .B(_22426_),
    .CO(_22427_),
    .S(_22428_));
 HA_X1 _41981_ (.A(\g_reduce0[12].adder.x[13] ),
    .B(_22429_),
    .CO(_22430_),
    .S(_22431_));
 HA_X1 _41982_ (.A(\g_reduce0[12].adder.x[12] ),
    .B(_22432_),
    .CO(_22433_),
    .S(_22434_));
 HA_X1 _41983_ (.A(\g_reduce0[12].adder.x[11] ),
    .B(_22435_),
    .CO(_22436_),
    .S(_22437_));
 HA_X1 _41984_ (.A(\g_reduce0[12].adder.x[9] ),
    .B(_22438_),
    .CO(_22439_),
    .S(_22440_));
 HA_X1 _41985_ (.A(\g_reduce0[12].adder.x[8] ),
    .B(_22441_),
    .CO(_22442_),
    .S(_22443_));
 HA_X1 _41986_ (.A(\g_reduce0[12].adder.x[7] ),
    .B(_22444_),
    .CO(_22445_),
    .S(_22446_));
 HA_X1 _41987_ (.A(\g_reduce0[12].adder.x[6] ),
    .B(_22447_),
    .CO(_22448_),
    .S(_22449_));
 HA_X1 _41988_ (.A(\g_reduce0[12].adder.x[5] ),
    .B(_22450_),
    .CO(_22451_),
    .S(_22452_));
 HA_X1 _41989_ (.A(\g_reduce0[12].adder.x[4] ),
    .B(_22453_),
    .CO(_22454_),
    .S(_22455_));
 HA_X1 _41990_ (.A(\g_reduce0[12].adder.x[3] ),
    .B(_22456_),
    .CO(_22457_),
    .S(_22458_));
 HA_X1 _41991_ (.A(\g_reduce0[12].adder.x[2] ),
    .B(_22459_),
    .CO(_22460_),
    .S(_22461_));
 HA_X1 _41992_ (.A(\g_reduce0[12].adder.x[1] ),
    .B(_22462_),
    .CO(_22463_),
    .S(_22464_));
 HA_X1 _41993_ (.A(_22465_),
    .B(\g_reduce0[14].adder.x[0] ),
    .CO(_22466_),
    .S(_22467_));
 HA_X1 _41994_ (.A(_22468_),
    .B(\g_reduce0[14].adder.x[10] ),
    .CO(_22469_),
    .S(_22470_));
 HA_X1 _41995_ (.A(_22471_),
    .B(_22437_),
    .CO(_22472_),
    .S(_22473_));
 HA_X1 _41996_ (.A(\g_reduce0[12].adder.x[14] ),
    .B(_22474_),
    .CO(_22475_),
    .S(_22476_));
 HA_X1 _41997_ (.A(_14196_),
    .B(_14197_),
    .CO(_22477_),
    .S(_22478_));
 HA_X1 _41998_ (.A(_14196_),
    .B(_14201_),
    .CO(_22479_),
    .S(_22480_));
 HA_X1 _41999_ (.A(_22481_),
    .B(_22482_),
    .CO(_22483_),
    .S(_22484_));
 HA_X1 _42000_ (.A(_22485_),
    .B(_22486_),
    .CO(_22487_),
    .S(_22488_));
 HA_X1 _42001_ (.A(_22485_),
    .B(_22489_),
    .CO(_22490_),
    .S(_22491_));
 HA_X1 _42002_ (.A(_22492_),
    .B(_22493_),
    .CO(_22494_),
    .S(_22495_));
 HA_X1 _42003_ (.A(_22496_),
    .B(_22493_),
    .CO(_22497_),
    .S(_22498_));
 HA_X1 _42004_ (.A(_22499_),
    .B(_22500_),
    .CO(_22501_),
    .S(_22502_));
 HA_X1 _42005_ (.A(_22503_),
    .B(_22500_),
    .CO(_22504_),
    .S(_22505_));
 HA_X1 _42006_ (.A(_22506_),
    .B(_22507_),
    .CO(_22508_),
    .S(_22509_));
 HA_X1 _42007_ (.A(_22506_),
    .B(_22510_),
    .CO(_22511_),
    .S(_22512_));
 HA_X1 _42008_ (.A(_22513_),
    .B(_22514_),
    .CO(_22515_),
    .S(_22516_));
 HA_X1 _42009_ (.A(_22517_),
    .B(_22514_),
    .CO(_22518_),
    .S(_22519_));
 HA_X1 _42010_ (.A(_22520_),
    .B(_22521_),
    .CO(_22522_),
    .S(_22523_));
 HA_X1 _42011_ (.A(_22524_),
    .B(_22521_),
    .CO(_22525_),
    .S(_22526_));
 HA_X1 _42012_ (.A(_22482_),
    .B(_22527_),
    .CO(_22528_),
    .S(_22529_));
 HA_X1 _42013_ (.A(_22530_),
    .B(_22531_),
    .CO(_22532_),
    .S(_22533_));
 HA_X1 _42014_ (.A(_22530_),
    .B(_22534_),
    .CO(_22535_),
    .S(_22536_));
 HA_X1 _42015_ (.A(_22537_),
    .B(_22538_),
    .CO(_14195_),
    .S(_22539_));
 HA_X1 _42016_ (.A(_22537_),
    .B(_22540_),
    .CO(_14200_),
    .S(_22541_));
 HA_X1 _42017_ (.A(_22542_),
    .B(_22543_),
    .CO(_22544_),
    .S(_14209_));
 HA_X1 _42018_ (.A(_22545_),
    .B(_22543_),
    .CO(_22546_),
    .S(_22547_));
 HA_X1 _42019_ (.A(_22545_),
    .B(_22543_),
    .CO(_22548_),
    .S(_22549_));
 HA_X1 _42020_ (.A(_22550_),
    .B(_22551_),
    .CO(_22552_),
    .S(_22553_));
 HA_X1 _42021_ (.A(_22542_),
    .B(_22554_),
    .CO(_14206_),
    .S(_22555_));
 HA_X1 _42022_ (.A(_22556_),
    .B(_22557_),
    .CO(_19429_),
    .S(_22558_));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_0_clk));
 DFFR_X1 \g_reduce0[0].adder.x[0]$_DFF_PN0_  (.D(_00000_),
    .RN(net348),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[0].adder.x[0] ),
    .QN(_00562_));
 DFFR_X2 \g_reduce0[0].adder.x[10]$_DFF_PN0_  (.D(_00001_),
    .RN(net349),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[0].adder.x[10] ),
    .QN(_13268_));
 DFFR_X2 \g_reduce0[0].adder.x[11]$_DFF_PN0_  (.D(_00002_),
    .RN(net348),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[0].adder.x[11] ),
    .QN(_21997_));
 DFFR_X2 \g_reduce0[0].adder.x[12]$_DFF_PN0_  (.D(_00003_),
    .RN(net349),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[0].adder.x[12] ),
    .QN(_21994_));
 DFFR_X1 \g_reduce0[0].adder.x[13]$_DFF_PN0_  (.D(_00004_),
    .RN(net349),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[0].adder.x[13] ),
    .QN(_21991_));
 DFFR_X2 \g_reduce0[0].adder.x[14]$_DFF_PN0_  (.D(_00005_),
    .RN(net349),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[0].adder.x[14] ),
    .QN(_22033_));
 DFFR_X2 \g_reduce0[0].adder.x[15]$_DFF_PN0_  (.D(_00006_),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_reduce0[0].adder.x[15] ),
    .QN(_13269_));
 DFFR_X1 \g_reduce0[0].adder.x[1]$_DFF_PN0_  (.D(_00007_),
    .RN(net348),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[0].adder.x[1] ),
    .QN(_22027_));
 DFFR_X1 \g_reduce0[0].adder.x[2]$_DFF_PN0_  (.D(_00008_),
    .RN(net348),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[0].adder.x[2] ),
    .QN(_22024_));
 DFFR_X1 \g_reduce0[0].adder.x[3]$_DFF_PN0_  (.D(_00009_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[0].adder.x[3] ),
    .QN(_22021_));
 DFFR_X1 \g_reduce0[0].adder.x[4]$_DFF_PN0_  (.D(_00010_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[0].adder.x[4] ),
    .QN(_22018_));
 DFFR_X1 \g_reduce0[0].adder.x[5]$_DFF_PN0_  (.D(_00011_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[0].adder.x[5] ),
    .QN(_22015_));
 DFFR_X1 \g_reduce0[0].adder.x[6]$_DFF_PN0_  (.D(_00012_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[0].adder.x[6] ),
    .QN(_22012_));
 DFFR_X1 \g_reduce0[0].adder.x[7]$_DFF_PN0_  (.D(_00013_),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_reduce0[0].adder.x[7] ),
    .QN(_22009_));
 DFFR_X2 \g_reduce0[0].adder.x[8]$_DFF_PN0_  (.D(_00014_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[0].adder.x[8] ),
    .QN(_22006_));
 DFFR_X1 \g_reduce0[0].adder.x[9]$_DFF_PN0_  (.D(_00015_),
    .RN(net348),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[0].adder.x[9] ),
    .QN(_22003_));
 DFFR_X1 \g_reduce0[10].adder.x[0]$_DFF_PN0_  (.D(_00016_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.x[0] ),
    .QN(_00589_));
 DFFR_X1 \g_reduce0[10].adder.x[10]$_DFF_PN0_  (.D(_00017_),
    .RN(net347),
    .CK(clknet_leaf_74_clk),
    .Q(\g_reduce0[10].adder.x[10] ),
    .QN(_00590_));
 DFFR_X2 \g_reduce0[10].adder.x[11]$_DFF_PN0_  (.D(_00018_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[10].adder.x[11] ),
    .QN(_22288_));
 DFFR_X2 \g_reduce0[10].adder.x[12]$_DFF_PN0_  (.D(_00019_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.x[12] ),
    .QN(_22285_));
 DFFR_X1 \g_reduce0[10].adder.x[13]$_DFF_PN0_  (.D(_00020_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.x[13] ),
    .QN(_22282_));
 DFFR_X1 \g_reduce0[10].adder.x[14]$_DFF_PN0_  (.D(_00021_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.x[14] ),
    .QN(_22327_));
 DFFR_X2 \g_reduce0[10].adder.x[15]$_DFF_PN0_  (.D(_00022_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[10].adder.x[15] ),
    .QN(_13270_));
 DFFR_X2 \g_reduce0[10].adder.x[1]$_DFF_PN0_  (.D(_00023_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.x[1] ),
    .QN(_22315_));
 DFFR_X2 \g_reduce0[10].adder.x[2]$_DFF_PN0_  (.D(_00024_),
    .RN(net347),
    .CK(clknet_leaf_74_clk),
    .Q(\g_reduce0[10].adder.x[2] ),
    .QN(_22312_));
 DFFR_X2 \g_reduce0[10].adder.x[3]$_DFF_PN0_  (.D(_00025_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.x[3] ),
    .QN(_22309_));
 DFFR_X2 \g_reduce0[10].adder.x[4]$_DFF_PN0_  (.D(_00026_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.x[4] ),
    .QN(_22306_));
 DFFR_X2 \g_reduce0[10].adder.x[5]$_DFF_PN0_  (.D(_00027_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.x[5] ),
    .QN(_22303_));
 DFFR_X2 \g_reduce0[10].adder.x[6]$_DFF_PN0_  (.D(_00028_),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(\g_reduce0[10].adder.x[6] ),
    .QN(_22300_));
 DFFR_X2 \g_reduce0[10].adder.x[7]$_DFF_PN0_  (.D(_00029_),
    .RN(net347),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.x[7] ),
    .QN(_22297_));
 DFFR_X2 \g_reduce0[10].adder.x[8]$_DFF_PN0_  (.D(_00030_),
    .RN(net347),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.x[8] ),
    .QN(_22294_));
 DFFR_X2 \g_reduce0[10].adder.x[9]$_DFF_PN0_  (.D(_00031_),
    .RN(net346),
    .CK(clknet_leaf_74_clk),
    .Q(\g_reduce0[10].adder.x[9] ),
    .QN(_22291_));
 DFFR_X1 \g_reduce0[12].adder.x[0]$_DFF_PN0_  (.D(_00032_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[12].adder.x[0] ),
    .QN(_22465_));
 DFFR_X1 \g_reduce0[12].adder.x[10]$_DFF_PN0_  (.D(_00033_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[12].adder.x[10] ),
    .QN(_22468_));
 DFFR_X1 \g_reduce0[12].adder.x[11]$_DFF_PN0_  (.D(_00034_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[12].adder.x[11] ),
    .QN(_00607_));
 DFFR_X1 \g_reduce0[12].adder.x[12]$_DFF_PN0_  (.D(_00035_),
    .RN(net348),
    .CK(clknet_leaf_129_clk),
    .Q(\g_reduce0[12].adder.x[12] ),
    .QN(_00612_));
 DFFR_X1 \g_reduce0[12].adder.x[13]$_DFF_PN0_  (.D(_00036_),
    .RN(net348),
    .CK(clknet_leaf_129_clk),
    .Q(\g_reduce0[12].adder.x[13] ),
    .QN(_00615_));
 DFFR_X1 \g_reduce0[12].adder.x[14]$_DFF_PN0_  (.D(_00037_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[12].adder.x[14] ),
    .QN(_13271_));
 DFFR_X2 \g_reduce0[12].adder.x[15]$_DFF_PN0_  (.D(_00038_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[12].adder.x[15] ),
    .QN(_13272_));
 DFFR_X1 \g_reduce0[12].adder.x[1]$_DFF_PN0_  (.D(_00039_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[1] ),
    .QN(_00602_));
 DFFR_X1 \g_reduce0[12].adder.x[2]$_DFF_PN0_  (.D(_00040_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[2] ),
    .QN(_00606_));
 DFFR_X1 \g_reduce0[12].adder.x[3]$_DFF_PN0_  (.D(_00041_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[3] ),
    .QN(_00605_));
 DFFR_X1 \g_reduce0[12].adder.x[4]$_DFF_PN0_  (.D(_00042_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[4] ),
    .QN(_00609_));
 DFFR_X1 \g_reduce0[12].adder.x[5]$_DFF_PN0_  (.D(_00043_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[12].adder.x[5] ),
    .QN(_00608_));
 DFFR_X1 \g_reduce0[12].adder.x[6]$_DFF_PN0_  (.D(_00044_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[12].adder.x[6] ),
    .QN(_00611_));
 DFFR_X2 \g_reduce0[12].adder.x[7]$_DFF_PN0_  (.D(_00045_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[12].adder.x[7] ),
    .QN(_00610_));
 DFFR_X2 \g_reduce0[12].adder.x[8]$_DFF_PN0_  (.D(_00046_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[8] ),
    .QN(_00614_));
 DFFR_X1 \g_reduce0[12].adder.x[9]$_DFF_PN0_  (.D(_00047_),
    .RN(net348),
    .CK(clknet_leaf_118_clk),
    .Q(\g_reduce0[12].adder.x[9] ),
    .QN(_00613_));
 DFFR_X1 \g_reduce0[14].adder.x[0]$_DFF_PN0_  (.D(_00048_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[14].adder.x[0] ),
    .QN(_00603_));
 DFFR_X1 \g_reduce0[14].adder.x[10]$_DFF_PN0_  (.D(_00049_),
    .RN(net348),
    .CK(clknet_leaf_127_clk),
    .Q(\g_reduce0[14].adder.x[10] ),
    .QN(_00604_));
 DFFR_X2 \g_reduce0[14].adder.x[11]$_DFF_PN0_  (.D(_00050_),
    .RN(net348),
    .CK(clknet_leaf_126_clk),
    .Q(\g_reduce0[14].adder.x[11] ),
    .QN(_22435_));
 DFFR_X2 \g_reduce0[14].adder.x[12]$_DFF_PN0_  (.D(_00051_),
    .RN(net348),
    .CK(clknet_leaf_126_clk),
    .Q(\g_reduce0[14].adder.x[12] ),
    .QN(_22432_));
 DFFR_X1 \g_reduce0[14].adder.x[13]$_DFF_PN0_  (.D(_00052_),
    .RN(net348),
    .CK(clknet_leaf_129_clk),
    .Q(\g_reduce0[14].adder.x[13] ),
    .QN(_22429_));
 DFFR_X1 \g_reduce0[14].adder.x[14]$_DFF_PN0_  (.D(_00053_),
    .RN(net348),
    .CK(clknet_leaf_129_clk),
    .Q(\g_reduce0[14].adder.x[14] ),
    .QN(_22474_));
 DFFR_X2 \g_reduce0[14].adder.x[15]$_DFF_PN0_  (.D(_00054_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[14].adder.x[15] ),
    .QN(_13273_));
 DFFR_X1 \g_reduce0[14].adder.x[1]$_DFF_PN0_  (.D(_00055_),
    .RN(net348),
    .CK(clknet_leaf_126_clk),
    .Q(\g_reduce0[14].adder.x[1] ),
    .QN(_22462_));
 DFFR_X2 \g_reduce0[14].adder.x[2]$_DFF_PN0_  (.D(_00056_),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_reduce0[14].adder.x[2] ),
    .QN(_22459_));
 DFFR_X1 \g_reduce0[14].adder.x[3]$_DFF_PN0_  (.D(_00057_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[14].adder.x[3] ),
    .QN(_22456_));
 DFFR_X1 \g_reduce0[14].adder.x[4]$_DFF_PN0_  (.D(_00058_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[14].adder.x[4] ),
    .QN(_22453_));
 DFFR_X1 \g_reduce0[14].adder.x[5]$_DFF_PN0_  (.D(_00059_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[14].adder.x[5] ),
    .QN(_22450_));
 DFFR_X1 \g_reduce0[14].adder.x[6]$_DFF_PN0_  (.D(_00060_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[14].adder.x[6] ),
    .QN(_22447_));
 DFFR_X1 \g_reduce0[14].adder.x[7]$_DFF_PN0_  (.D(_00061_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.x[7] ),
    .QN(_22444_));
 DFFR_X1 \g_reduce0[14].adder.x[8]$_DFF_PN0_  (.D(_00062_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.x[8] ),
    .QN(_22441_));
 DFFR_X1 \g_reduce0[14].adder.x[9]$_DFF_PN0_  (.D(_00063_),
    .RN(net348),
    .CK(clknet_leaf_119_clk),
    .Q(\g_reduce0[14].adder.x[9] ),
    .QN(_22438_));
 DFFR_X1 \g_reduce0[2].adder.x[0]$_DFF_PN0_  (.D(_00064_),
    .RN(net348),
    .CK(clknet_leaf_130_clk),
    .Q(\g_reduce0[2].adder.x[0] ),
    .QN(_00561_));
 DFFR_X1 \g_reduce0[2].adder.x[10]$_DFF_PN0_  (.D(_00065_),
    .RN(net348),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[2].adder.x[10] ),
    .QN(_22000_));
 DFFR_X1 \g_reduce0[2].adder.x[11]$_DFF_PN0_  (.D(_00066_),
    .RN(net348),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[2].adder.x[11] ),
    .QN(_00565_));
 DFFR_X2 \g_reduce0[2].adder.x[12]$_DFF_PN0_  (.D(_00067_),
    .RN(net349),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[2].adder.x[12] ),
    .QN(_00570_));
 DFFR_X1 \g_reduce0[2].adder.x[13]$_DFF_PN0_  (.D(_00068_),
    .RN(net349),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[2].adder.x[13] ),
    .QN(_00573_));
 DFFR_X2 \g_reduce0[2].adder.x[14]$_DFF_PN0_  (.D(_00069_),
    .RN(net348),
    .CK(clknet_leaf_135_clk),
    .Q(\g_reduce0[2].adder.x[14] ),
    .QN(_13274_));
 DFFR_X1 \g_reduce0[2].adder.x[15]$_DFF_PN0_  (.D(_00070_),
    .RN(net348),
    .CK(clknet_leaf_130_clk),
    .Q(\g_reduce0[2].adder.x[15] ),
    .QN(_13275_));
 DFFR_X1 \g_reduce0[2].adder.x[1]$_DFF_PN0_  (.D(_00071_),
    .RN(net348),
    .CK(clknet_leaf_129_clk),
    .Q(\g_reduce0[2].adder.x[1] ),
    .QN(_00560_));
 DFFR_X1 \g_reduce0[2].adder.x[2]$_DFF_PN0_  (.D(_00072_),
    .RN(net348),
    .CK(clknet_leaf_139_clk),
    .Q(\g_reduce0[2].adder.x[2] ),
    .QN(_00564_));
 DFFR_X1 \g_reduce0[2].adder.x[3]$_DFF_PN0_  (.D(_00073_),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_reduce0[2].adder.x[3] ),
    .QN(_00563_));
 DFFR_X1 \g_reduce0[2].adder.x[4]$_DFF_PN0_  (.D(_00074_),
    .RN(net348),
    .CK(clknet_leaf_136_clk),
    .Q(\g_reduce0[2].adder.x[4] ),
    .QN(_00567_));
 DFFR_X1 \g_reduce0[2].adder.x[5]$_DFF_PN0_  (.D(_00075_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[2].adder.x[5] ),
    .QN(_00566_));
 DFFR_X1 \g_reduce0[2].adder.x[6]$_DFF_PN0_  (.D(_00076_),
    .RN(net348),
    .CK(clknet_leaf_130_clk),
    .Q(\g_reduce0[2].adder.x[6] ),
    .QN(_00569_));
 DFFR_X1 \g_reduce0[2].adder.x[7]$_DFF_PN0_  (.D(_00077_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[2].adder.x[7] ),
    .QN(_00568_));
 DFFR_X1 \g_reduce0[2].adder.x[8]$_DFF_PN0_  (.D(_00078_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[2].adder.x[8] ),
    .QN(_00572_));
 DFFR_X1 \g_reduce0[2].adder.x[9]$_DFF_PN0_  (.D(_00079_),
    .RN(net348),
    .CK(clknet_leaf_137_clk),
    .Q(\g_reduce0[2].adder.x[9] ),
    .QN(_00571_));
 DFFR_X1 \g_reduce0[4].adder.x[0]$_DFF_PN0_  (.D(_00080_),
    .RN(net349),
    .CK(clknet_leaf_111_clk),
    .Q(\g_reduce0[4].adder.x[0] ),
    .QN(_22171_));
 DFFR_X2 \g_reduce0[4].adder.x[10]$_DFF_PN0_  (.D(_00081_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[4].adder.x[10] ),
    .QN(_22174_));
 DFFR_X1 \g_reduce0[4].adder.x[11]$_DFF_PN0_  (.D(_00082_),
    .RN(net346),
    .CK(clknet_leaf_104_clk),
    .Q(\g_reduce0[4].adder.x[11] ),
    .QN(_00579_));
 DFFR_X1 \g_reduce0[4].adder.x[12]$_DFF_PN0_  (.D(_00083_),
    .RN(net346),
    .CK(clknet_leaf_104_clk),
    .Q(\g_reduce0[4].adder.x[12] ),
    .QN(_00584_));
 DFFR_X1 \g_reduce0[4].adder.x[13]$_DFF_PN0_  (.D(_00084_),
    .RN(net346),
    .CK(clknet_leaf_104_clk),
    .Q(\g_reduce0[4].adder.x[13] ),
    .QN(_00587_));
 DFFR_X2 \g_reduce0[4].adder.x[14]$_DFF_PN0_  (.D(_00085_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[4].adder.x[14] ),
    .QN(_13276_));
 DFFR_X2 \g_reduce0[4].adder.x[15]$_DFF_PN0_  (.D(_00086_),
    .RN(net349),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[4].adder.x[15] ),
    .QN(_13277_));
 DFFR_X1 \g_reduce0[4].adder.x[1]$_DFF_PN0_  (.D(_00087_),
    .RN(net349),
    .CK(clknet_leaf_111_clk),
    .Q(\g_reduce0[4].adder.x[1] ),
    .QN(_00574_));
 DFFR_X1 \g_reduce0[4].adder.x[2]$_DFF_PN0_  (.D(_00088_),
    .RN(net349),
    .CK(clknet_leaf_111_clk),
    .Q(\g_reduce0[4].adder.x[2] ),
    .QN(_00578_));
 DFFR_X2 \g_reduce0[4].adder.x[3]$_DFF_PN0_  (.D(_00089_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[4].adder.x[3] ),
    .QN(_00577_));
 DFFR_X1 \g_reduce0[4].adder.x[4]$_DFF_PN0_  (.D(_00090_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[4].adder.x[4] ),
    .QN(_00581_));
 DFFR_X2 \g_reduce0[4].adder.x[5]$_DFF_PN0_  (.D(_00091_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[4].adder.x[5] ),
    .QN(_00580_));
 DFFR_X2 \g_reduce0[4].adder.x[6]$_DFF_PN0_  (.D(_00092_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[4].adder.x[6] ),
    .QN(_00583_));
 DFFR_X2 \g_reduce0[4].adder.x[7]$_DFF_PN0_  (.D(_00093_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[4].adder.x[7] ),
    .QN(_00582_));
 DFFR_X2 \g_reduce0[4].adder.x[8]$_DFF_PN0_  (.D(_00094_),
    .RN(net349),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[4].adder.x[8] ),
    .QN(_00586_));
 DFFR_X2 \g_reduce0[4].adder.x[9]$_DFF_PN0_  (.D(_00095_),
    .RN(net349),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[4].adder.x[9] ),
    .QN(_00585_));
 DFFR_X1 \g_reduce0[6].adder.x[0]$_DFF_PN0_  (.D(_00096_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[0] ),
    .QN(_00575_));
 DFFR_X1 \g_reduce0[6].adder.x[10]$_DFF_PN0_  (.D(_00097_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[10] ),
    .QN(_00576_));
 DFFR_X1 \g_reduce0[6].adder.x[11]$_DFF_PN0_  (.D(_00098_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[11] ),
    .QN(_22141_));
 DFFR_X1 \g_reduce0[6].adder.x[12]$_DFF_PN0_  (.D(_00099_),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(\g_reduce0[6].adder.x[12] ),
    .QN(_22138_));
 DFFR_X1 \g_reduce0[6].adder.x[13]$_DFF_PN0_  (.D(_00100_),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(\g_reduce0[6].adder.x[13] ),
    .QN(_22135_));
 DFFR_X1 \g_reduce0[6].adder.x[14]$_DFF_PN0_  (.D(_00101_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[14] ),
    .QN(_22180_));
 DFFR_X2 \g_reduce0[6].adder.x[15]$_DFF_PN0_  (.D(_00102_),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(\g_reduce0[6].adder.x[15] ),
    .QN(_13278_));
 DFFR_X2 \g_reduce0[6].adder.x[1]$_DFF_PN0_  (.D(_00103_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[1] ),
    .QN(_22168_));
 DFFR_X1 \g_reduce0[6].adder.x[2]$_DFF_PN0_  (.D(_00104_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[2] ),
    .QN(_22165_));
 DFFR_X2 \g_reduce0[6].adder.x[3]$_DFF_PN0_  (.D(_00105_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[3] ),
    .QN(_22162_));
 DFFR_X1 \g_reduce0[6].adder.x[4]$_DFF_PN0_  (.D(_00106_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[4] ),
    .QN(_22159_));
 DFFR_X2 \g_reduce0[6].adder.x[5]$_DFF_PN0_  (.D(_00107_),
    .RN(net346),
    .CK(clknet_leaf_104_clk),
    .Q(\g_reduce0[6].adder.x[5] ),
    .QN(_22156_));
 DFFR_X2 \g_reduce0[6].adder.x[6]$_DFF_PN0_  (.D(_00108_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[6] ),
    .QN(_22153_));
 DFFR_X2 \g_reduce0[6].adder.x[7]$_DFF_PN0_  (.D(_00109_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[7] ),
    .QN(_22150_));
 DFFR_X2 \g_reduce0[6].adder.x[8]$_DFF_PN0_  (.D(_00110_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.x[8] ),
    .QN(_22147_));
 DFFR_X2 \g_reduce0[6].adder.x[9]$_DFF_PN0_  (.D(_00111_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.x[9] ),
    .QN(_22144_));
 DFFR_X1 \g_reduce0[8].adder.x[0]$_DFF_PN0_  (.D(_00112_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[0] ),
    .QN(_22318_));
 DFFR_X1 \g_reduce0[8].adder.x[10]$_DFF_PN0_  (.D(_00113_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[10] ),
    .QN(_22321_));
 DFFR_X1 \g_reduce0[8].adder.x[11]$_DFF_PN0_  (.D(_00114_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[8].adder.x[11] ),
    .QN(_00593_));
 DFFR_X1 \g_reduce0[8].adder.x[12]$_DFF_PN0_  (.D(_00115_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[8].adder.x[12] ),
    .QN(_00598_));
 DFFR_X2 \g_reduce0[8].adder.x[13]$_DFF_PN0_  (.D(_00116_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[8].adder.x[13] ),
    .QN(_00601_));
 DFFR_X1 \g_reduce0[8].adder.x[14]$_DFF_PN0_  (.D(_00117_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[8].adder.x[14] ),
    .QN(_13279_));
 DFFR_X2 \g_reduce0[8].adder.x[15]$_DFF_PN0_  (.D(_00118_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[15] ),
    .QN(_13280_));
 DFFR_X1 \g_reduce0[8].adder.x[1]$_DFF_PN0_  (.D(_00119_),
    .RN(net347),
    .CK(clknet_leaf_70_clk),
    .Q(\g_reduce0[8].adder.x[1] ),
    .QN(_00588_));
 DFFR_X2 \g_reduce0[8].adder.x[2]$_DFF_PN0_  (.D(_00120_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[8].adder.x[2] ),
    .QN(_00592_));
 DFFR_X1 \g_reduce0[8].adder.x[3]$_DFF_PN0_  (.D(_00121_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[8].adder.x[3] ),
    .QN(_00591_));
 DFFR_X2 \g_reduce0[8].adder.x[4]$_DFF_PN0_  (.D(_00122_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[8].adder.x[4] ),
    .QN(_00595_));
 DFFR_X1 \g_reduce0[8].adder.x[5]$_DFF_PN0_  (.D(_00123_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[8].adder.x[5] ),
    .QN(_00594_));
 DFFR_X2 \g_reduce0[8].adder.x[6]$_DFF_PN0_  (.D(_00124_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[8].adder.x[6] ),
    .QN(_00597_));
 DFFR_X2 \g_reduce0[8].adder.x[7]$_DFF_PN0_  (.D(_00125_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[7] ),
    .QN(_00596_));
 DFFR_X1 \g_reduce0[8].adder.x[8]$_DFF_PN0_  (.D(_00126_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[8] ),
    .QN(_00600_));
 DFFR_X1 \g_reduce0[8].adder.x[9]$_DFF_PN0_  (.D(_00127_),
    .RN(net347),
    .CK(clknet_leaf_69_clk),
    .Q(\g_reduce0[8].adder.x[9] ),
    .QN(_00599_));
 DFFR_X1 \g_reduce1[0].adder.x[0]$_DFF_PN0_  (.D(_00128_),
    .RN(net348),
    .CK(clknet_leaf_131_clk),
    .Q(net277),
    .QN(_13281_));
 DFFR_X1 \g_reduce1[0].adder.x[10]$_DFF_PN0_  (.D(_00129_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net278),
    .QN(_13282_));
 DFFR_X1 \g_reduce1[0].adder.x[11]$_DFF_PN0_  (.D(_00130_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net279),
    .QN(_13283_));
 DFFR_X1 \g_reduce1[0].adder.x[12]$_DFF_PN0_  (.D(_00131_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net280),
    .QN(_13284_));
 DFFR_X1 \g_reduce1[0].adder.x[13]$_DFF_PN0_  (.D(_00132_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net281),
    .QN(_13285_));
 DFFR_X1 \g_reduce1[0].adder.x[14]$_DFF_PN0_  (.D(_00133_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net282),
    .QN(_13286_));
 DFFR_X1 \g_reduce1[0].adder.x[15]$_DFF_PN0_  (.D(_00134_),
    .RN(net348),
    .CK(clknet_leaf_131_clk),
    .Q(net283),
    .QN(_13287_));
 DFFR_X1 \g_reduce1[0].adder.x[1]$_DFF_PN0_  (.D(_00135_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net288),
    .QN(_13288_));
 DFFR_X1 \g_reduce1[0].adder.x[2]$_DFF_PN0_  (.D(_00136_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net299),
    .QN(_13289_));
 DFFR_X1 \g_reduce1[0].adder.x[3]$_DFF_PN0_  (.D(_00137_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net310),
    .QN(_13290_));
 DFFR_X1 \g_reduce1[0].adder.x[4]$_DFF_PN0_  (.D(_00138_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net321),
    .QN(_13291_));
 DFFR_X1 \g_reduce1[0].adder.x[5]$_DFF_PN0_  (.D(_00139_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net332),
    .QN(_13292_));
 DFFR_X1 \g_reduce1[0].adder.x[6]$_DFF_PN0_  (.D(_00140_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net337),
    .QN(_13293_));
 DFFR_X1 \g_reduce1[0].adder.x[7]$_DFF_PN0_  (.D(_00141_),
    .RN(net349),
    .CK(clknet_leaf_133_clk),
    .Q(net338),
    .QN(_13294_));
 DFFR_X1 \g_reduce1[0].adder.x[8]$_DFF_PN0_  (.D(_00142_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net339),
    .QN(_13295_));
 DFFR_X1 \g_reduce1[0].adder.x[9]$_DFF_PN0_  (.D(_00143_),
    .RN(net349),
    .CK(clknet_leaf_132_clk),
    .Q(net340),
    .QN(_13296_));
 DFFR_X1 \g_reduce1[2].adder.x[0]$_DFF_PN0_  (.D(_00144_),
    .RN(net346),
    .CK(clknet_leaf_100_clk),
    .Q(net284),
    .QN(_13297_));
 DFFR_X1 \g_reduce1[2].adder.x[10]$_DFF_PN0_  (.D(_00145_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net295),
    .QN(_13298_));
 DFFR_X1 \g_reduce1[2].adder.x[11]$_DFF_PN0_  (.D(_00146_),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(net296),
    .QN(_13299_));
 DFFR_X1 \g_reduce1[2].adder.x[12]$_DFF_PN0_  (.D(_00147_),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(net297),
    .QN(_13300_));
 DFFR_X1 \g_reduce1[2].adder.x[13]$_DFF_PN0_  (.D(_00148_),
    .RN(net346),
    .CK(clknet_leaf_100_clk),
    .Q(net298),
    .QN(_13301_));
 DFFR_X1 \g_reduce1[2].adder.x[14]$_DFF_PN0_  (.D(_00149_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net300),
    .QN(_13302_));
 DFFR_X1 \g_reduce1[2].adder.x[15]$_DFF_PN0_  (.D(_00150_),
    .RN(net346),
    .CK(clknet_leaf_100_clk),
    .Q(net301),
    .QN(_13303_));
 DFFR_X1 \g_reduce1[2].adder.x[1]$_DFF_PN0_  (.D(_00151_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net285),
    .QN(_13304_));
 DFFR_X1 \g_reduce1[2].adder.x[2]$_DFF_PN0_  (.D(_00152_),
    .RN(net346),
    .CK(clknet_leaf_98_clk),
    .Q(net286),
    .QN(_13305_));
 DFFR_X1 \g_reduce1[2].adder.x[3]$_DFF_PN0_  (.D(_00153_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net287),
    .QN(_13306_));
 DFFR_X1 \g_reduce1[2].adder.x[4]$_DFF_PN0_  (.D(_00154_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net289),
    .QN(_13307_));
 DFFR_X1 \g_reduce1[2].adder.x[5]$_DFF_PN0_  (.D(_00155_),
    .RN(net346),
    .CK(clknet_leaf_98_clk),
    .Q(net290),
    .QN(_13308_));
 DFFR_X1 \g_reduce1[2].adder.x[6]$_DFF_PN0_  (.D(_00156_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net291),
    .QN(_13309_));
 DFFR_X1 \g_reduce1[2].adder.x[7]$_DFF_PN0_  (.D(_00157_),
    .RN(net346),
    .CK(clknet_leaf_100_clk),
    .Q(net292),
    .QN(_13310_));
 DFFR_X1 \g_reduce1[2].adder.x[8]$_DFF_PN0_  (.D(_00158_),
    .RN(net346),
    .CK(clknet_leaf_98_clk),
    .Q(net293),
    .QN(_13311_));
 DFFR_X1 \g_reduce1[2].adder.x[9]$_DFF_PN0_  (.D(_00159_),
    .RN(net346),
    .CK(clknet_leaf_99_clk),
    .Q(net294),
    .QN(_13312_));
 DFFR_X1 \g_reduce1[4].adder.x[0]$_DFF_PN0_  (.D(_00160_),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(net302),
    .QN(_13313_));
 DFFR_X1 \g_reduce1[4].adder.x[10]$_DFF_PN0_  (.D(_00161_),
    .RN(net346),
    .CK(clknet_leaf_77_clk),
    .Q(net313),
    .QN(_13314_));
 DFFR_X1 \g_reduce1[4].adder.x[11]$_DFF_PN0_  (.D(_00162_),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(net314),
    .QN(_13315_));
 DFFR_X2 \g_reduce1[4].adder.x[12]$_DFF_PN0_  (.D(_00163_),
    .RN(net347),
    .CK(clknet_leaf_74_clk),
    .Q(net315),
    .QN(_13316_));
 DFFR_X2 \g_reduce1[4].adder.x[13]$_DFF_PN0_  (.D(_00164_),
    .RN(net346),
    .CK(clknet_leaf_74_clk),
    .Q(net316),
    .QN(_13317_));
 DFFR_X2 \g_reduce1[4].adder.x[14]$_DFF_PN0_  (.D(_00165_),
    .RN(net347),
    .CK(clknet_leaf_74_clk),
    .Q(net317),
    .QN(_13318_));
 DFFR_X1 \g_reduce1[4].adder.x[15]$_DFF_PN0_  (.D(_00166_),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(net318),
    .QN(_13319_));
 DFFR_X1 \g_reduce1[4].adder.x[1]$_DFF_PN0_  (.D(_00167_),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(net303),
    .QN(_13320_));
 DFFR_X1 \g_reduce1[4].adder.x[2]$_DFF_PN0_  (.D(_00168_),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(net304),
    .QN(_13321_));
 DFFR_X1 \g_reduce1[4].adder.x[3]$_DFF_PN0_  (.D(_00169_),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(net305),
    .QN(_13322_));
 DFFR_X1 \g_reduce1[4].adder.x[4]$_DFF_PN0_  (.D(_00170_),
    .RN(net348),
    .CK(clknet_leaf_105_clk),
    .Q(net306),
    .QN(_13323_));
 DFFR_X1 \g_reduce1[4].adder.x[5]$_DFF_PN0_  (.D(_00171_),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(net307),
    .QN(_13324_));
 DFFR_X1 \g_reduce1[4].adder.x[6]$_DFF_PN0_  (.D(_00172_),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(net308),
    .QN(_13325_));
 DFFR_X2 \g_reduce1[4].adder.x[7]$_DFF_PN0_  (.D(_00173_),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(net309),
    .QN(_13326_));
 DFFR_X1 \g_reduce1[4].adder.x[8]$_DFF_PN0_  (.D(_00174_),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(net311),
    .QN(_13327_));
 DFFR_X1 \g_reduce1[4].adder.x[9]$_DFF_PN0_  (.D(_00175_),
    .RN(net348),
    .CK(clknet_leaf_105_clk),
    .Q(net312),
    .QN(_13328_));
 DFFR_X1 \g_reduce1[6].adder.x[0]$_DFF_PN0_  (.D(_00176_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net319),
    .QN(_13329_));
 DFFR_X1 \g_reduce1[6].adder.x[10]$_DFF_PN0_  (.D(_00177_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net330),
    .QN(_13330_));
 DFFR_X1 \g_reduce1[6].adder.x[11]$_DFF_PN0_  (.D(_00178_),
    .RN(net348),
    .CK(clknet_leaf_131_clk),
    .Q(net331),
    .QN(_13331_));
 DFFR_X1 \g_reduce1[6].adder.x[12]$_DFF_PN0_  (.D(_00179_),
    .RN(net348),
    .CK(clknet_leaf_126_clk),
    .Q(net333),
    .QN(_13332_));
 DFFR_X1 \g_reduce1[6].adder.x[13]$_DFF_PN0_  (.D(_00180_),
    .RN(net348),
    .CK(clknet_leaf_131_clk),
    .Q(net334),
    .QN(_13333_));
 DFFR_X1 \g_reduce1[6].adder.x[14]$_DFF_PN0_  (.D(_00181_),
    .RN(net348),
    .CK(clknet_leaf_130_clk),
    .Q(net335),
    .QN(_13334_));
 DFFR_X1 \g_reduce1[6].adder.x[15]$_DFF_PN0_  (.D(_00182_),
    .RN(net348),
    .CK(clknet_leaf_124_clk),
    .Q(net336),
    .QN(_13335_));
 DFFR_X1 \g_reduce1[6].adder.x[1]$_DFF_PN0_  (.D(_00183_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net320),
    .QN(_13336_));
 DFFR_X1 \g_reduce1[6].adder.x[2]$_DFF_PN0_  (.D(_00184_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net322),
    .QN(_13337_));
 DFFR_X1 \g_reduce1[6].adder.x[3]$_DFF_PN0_  (.D(_00185_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net323),
    .QN(_13338_));
 DFFR_X1 \g_reduce1[6].adder.x[4]$_DFF_PN0_  (.D(_00186_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net324),
    .QN(_13339_));
 DFFR_X1 \g_reduce1[6].adder.x[5]$_DFF_PN0_  (.D(_00187_),
    .RN(net348),
    .CK(clknet_leaf_126_clk),
    .Q(net325),
    .QN(_13340_));
 DFFR_X1 \g_reduce1[6].adder.x[6]$_DFF_PN0_  (.D(_00188_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net326),
    .QN(_13341_));
 DFFR_X1 \g_reduce1[6].adder.x[7]$_DFF_PN0_  (.D(_00189_),
    .RN(net348),
    .CK(clknet_leaf_131_clk),
    .Q(net327),
    .QN(_13342_));
 DFFR_X1 \g_reduce1[6].adder.x[8]$_DFF_PN0_  (.D(_00190_),
    .RN(net348),
    .CK(clknet_leaf_125_clk),
    .Q(net328),
    .QN(_13343_));
 DFFR_X1 \g_reduce1[6].adder.x[9]$_DFF_PN0_  (.D(_00191_),
    .RN(net348),
    .CK(clknet_leaf_124_clk),
    .Q(net329),
    .QN(_13344_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.expa[0]$_DFF_PN0_  (.D(net10),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14217_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expa[1]$_DFF_PN0_  (.D(net20),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14223_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expa[2]$_DFF_PN0_  (.D(net30),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13345_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expa[3]$_DFF_PN0_  (.D(net39),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13346_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.expa[4]$_DFF_PN0_  (.D(net50),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13347_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expb[0]$_DFF_PN0_  (.D(net233),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[0].fa.b ),
    .QN(_14216_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expb[1]$_DFF_PN0_  (.D(net234),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[1].fa.b ),
    .QN(_14222_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expb[2]$_DFF_PN0_  (.D(net235),
    .RN(net347),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[2].fa.b ),
    .QN(_13348_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.expb[3]$_DFF_PN0_  (.D(net236),
    .RN(net347),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[3].fa.b ),
    .QN(_13349_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.expb[4]$_DFF_PN0_  (.D(net237),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[0].g_col[0].mult.expAdder.g_intermediate[4].fa.b ),
    .QN(_13350_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.sign$_DFF_PN0_  (.D(_00207_),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_row[0].g_col[0].mult.sign ),
    .QN(_13351_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[0] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[0] ),
    .QN(_13352_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[10] ),
    .RN(net345),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[10] ),
    .QN(_13353_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[11] ),
    .RN(net351),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[11] ),
    .QN(_13354_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[12] ),
    .RN(net345),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[12] ),
    .QN(_13355_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[13] ),
    .RN(net351),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[13] ),
    .QN(_13356_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[14] ),
    .RN(net351),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[14] ),
    .QN(_13357_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[15] ),
    .RN(net351),
    .CK(clknet_leaf_37_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[15] ),
    .QN(_13358_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[16] ),
    .RN(net351),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[16] ),
    .QN(_13359_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[17] ),
    .RN(net351),
    .CK(clknet_leaf_38_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[17] ),
    .QN(_13360_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[18] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[18] ),
    .QN(_13361_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[19] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[19] ),
    .QN(_13362_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[1] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[1] ),
    .QN(_13363_));
 DFFR_X2 \g_row[0].g_col[0].mult.stage1.t1[20]$_DFF_PN0_  (.D(net354),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[20] ),
    .QN(_13364_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[2] ),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[2] ),
    .QN(_14211_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[3] ),
    .RN(net351),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[3] ),
    .QN(_13365_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[4] ),
    .RN(net351),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[4] ),
    .QN(_13366_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[5] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[5] ),
    .QN(_13367_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[6] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[6] ),
    .QN(_13368_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[7] ),
    .RN(net351),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[7] ),
    .QN(_13369_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[8] ),
    .RN(net351),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[8] ),
    .QN(_13370_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t1[9] ),
    .RN(net345),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.a[9] ),
    .QN(_13371_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[10] ),
    .RN(net351),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[10] ),
    .QN(_13372_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[11] ),
    .RN(net351),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[11] ),
    .QN(_13373_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[12] ),
    .RN(net351),
    .CK(clknet_leaf_40_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[12] ),
    .QN(_13374_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[13] ),
    .RN(net345),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[13] ),
    .QN(_13375_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[14] ),
    .RN(net351),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[14] ),
    .QN(_13376_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[15] ),
    .RN(net351),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[15] ),
    .QN(_13377_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[16] ),
    .RN(net351),
    .CK(clknet_leaf_37_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[16] ),
    .QN(_13378_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[17] ),
    .RN(net351),
    .CK(clknet_leaf_38_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[17] ),
    .QN(_13379_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[18] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[18] ),
    .QN(_13380_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[19] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[19] ),
    .QN(_13381_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[1] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[1] ),
    .QN(_13382_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[20] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[20] ),
    .QN(_13383_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[2] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[2] ),
    .QN(_14212_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[3] ),
    .RN(net351),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[3] ),
    .QN(_13384_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[4] ),
    .RN(net351),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[4] ),
    .QN(_13385_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[5] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[5] ),
    .QN(_13386_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[6] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[6] ),
    .QN(_13387_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[7] ),
    .RN(net351),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[7] ),
    .QN(_13388_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[8] ),
    .RN(net351),
    .CK(clknet_leaf_43_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[8] ),
    .QN(_13389_));
 DFFR_X1 \g_row[0].g_col[0].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.stage1.dadda.t2[9] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[0].g_col[0].mult.adder.b[9] ),
    .QN(_13390_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[0]$_DFF_PN0_  (.D(_00192_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[0] ),
    .QN(_20389_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[10]$_DFF_PN0_  (.D(_00193_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.a[10] ),
    .QN(_20392_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[11]$_DFF_PN0_  (.D(_00194_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.a[11] ),
    .QN(_00453_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[12]$_DFF_PN0_  (.D(_00195_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.a[12] ),
    .QN(_00458_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[13]$_DFF_PN0_  (.D(_00196_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.a[13] ),
    .QN(_00461_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[14]$_DFF_PN0_  (.D(_00197_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.a[14] ),
    .QN(_13391_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[15]$_DFF_PN0_  (.D(\g_row[0].g_col[0].mult.sign ),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_reduce0[0].adder.a[15] ),
    .QN(_13392_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[1]$_DFF_PN0_  (.D(_00198_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[1] ),
    .QN(_00448_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[2]$_DFF_PN0_  (.D(_00199_),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_reduce0[0].adder.a[2] ),
    .QN(_00452_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[3]$_DFF_PN0_  (.D(_00200_),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_reduce0[0].adder.a[3] ),
    .QN(_00451_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[4]$_DFF_PN0_  (.D(_00201_),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_reduce0[0].adder.a[4] ),
    .QN(_00455_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[5]$_DFF_PN0_  (.D(_00202_),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_reduce0[0].adder.a[5] ),
    .QN(_00454_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[6]$_DFF_PN0_  (.D(_00203_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[6] ),
    .QN(_00457_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[7]$_DFF_PN0_  (.D(_00204_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[7] ),
    .QN(_00456_));
 DFFR_X2 \g_row[0].g_col[0].mult.x[8]$_DFF_PN0_  (.D(_00205_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[8] ),
    .QN(_00460_));
 DFFR_X1 \g_row[0].g_col[0].mult.x[9]$_DFF_PN0_  (.D(_00206_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.a[9] ),
    .QN(_00459_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.expa[0]$_DFF_PN0_  (.D(net156),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14236_));
 DFFR_X2 \g_row[0].g_col[1].mult.stage1.expa[1]$_DFF_PN0_  (.D(net157),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14242_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.expa[2]$_DFF_PN0_  (.D(net158),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13393_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.expa[3]$_DFF_PN0_  (.D(net159),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13394_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.expa[4]$_DFF_PN0_  (.D(net161),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13395_));
 DFFR_X2 \g_row[0].g_col[1].mult.stage1.expb[0]$_DFF_PN0_  (.D(net244),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[0].fa.b ),
    .QN(_14235_));
 DFFR_X2 \g_row[0].g_col[1].mult.stage1.expb[1]$_DFF_PN0_  (.D(net245),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[1].fa.b ),
    .QN(_14241_));
 DFFR_X2 \g_row[0].g_col[1].mult.stage1.expb[2]$_DFF_PN0_  (.D(net246),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[2].fa.b ),
    .QN(_13396_));
 DFFR_X2 \g_row[0].g_col[1].mult.stage1.expb[3]$_DFF_PN0_  (.D(net247),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[3].fa.b ),
    .QN(_13397_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.expb[4]$_DFF_PN0_  (.D(net249),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[0].g_col[1].mult.expAdder.g_intermediate[4].fa.b ),
    .QN(_13398_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.sign$_DFF_PN0_  (.D(_00223_),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_row[0].g_col[1].mult.sign ),
    .QN(_13399_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[0] ),
    .RN(net350),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[0] ),
    .QN(_13400_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[10] ),
    .RN(net276),
    .CK(clknet_leaf_181_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[10] ),
    .QN(_13401_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[11] ),
    .RN(net276),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[11] ),
    .QN(_13402_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[12] ),
    .RN(net351),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[12] ),
    .QN(_13403_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[13] ),
    .RN(net351),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[13] ),
    .QN(_13404_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[14] ),
    .RN(net276),
    .CK(clknet_leaf_181_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[14] ),
    .QN(_13405_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[15] ),
    .RN(net276),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[15] ),
    .QN(_13406_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[16] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[16] ),
    .QN(_13407_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[17] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[17] ),
    .QN(_13408_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[18] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[18] ),
    .QN(_13409_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[19] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[19] ),
    .QN(_13410_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[1] ),
    .RN(net350),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[1] ),
    .QN(_13411_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[2] ),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[2] ),
    .QN(_14230_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[3] ),
    .RN(net350),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[3] ),
    .QN(_13412_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[4] ),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[4] ),
    .QN(_13413_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[5] ),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[5] ),
    .QN(_13414_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[6] ),
    .RN(net350),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[6] ),
    .QN(_13415_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[7] ),
    .RN(net276),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[7] ),
    .QN(_13416_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[8] ),
    .RN(net276),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[8] ),
    .QN(_13417_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t1[9] ),
    .RN(net276),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.a[9] ),
    .QN(_13418_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[10] ),
    .RN(net276),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[10] ),
    .QN(_13419_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[11] ),
    .RN(net276),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[11] ),
    .QN(_13420_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[12] ),
    .RN(net351),
    .CK(clknet_leaf_182_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[12] ),
    .QN(_13421_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[13] ),
    .RN(net276),
    .CK(clknet_leaf_181_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[13] ),
    .QN(_13422_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[14] ),
    .RN(net276),
    .CK(clknet_leaf_181_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[14] ),
    .QN(_13423_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[15] ),
    .RN(net276),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[15] ),
    .QN(_13424_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[16] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[16] ),
    .QN(_13425_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[17] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[17] ),
    .QN(_13426_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[18] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[18] ),
    .QN(_13427_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[19] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[19] ),
    .QN(_13428_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[1] ),
    .RN(net350),
    .CK(clknet_leaf_178_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[1] ),
    .QN(_13429_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[20] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[20] ),
    .QN(_13430_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[2] ),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[2] ),
    .QN(_14231_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[3] ),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[3] ),
    .QN(_13431_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[4] ),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[4] ),
    .QN(_13432_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[5] ),
    .RN(net350),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[5] ),
    .QN(_13433_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[6] ),
    .RN(net350),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[6] ),
    .QN(_13434_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[7] ),
    .RN(net276),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[7] ),
    .QN(_13435_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[8] ),
    .RN(net276),
    .CK(clknet_leaf_180_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[8] ),
    .QN(_13436_));
 DFFR_X1 \g_row[0].g_col[1].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.stage1.dadda.t2[9] ),
    .RN(net276),
    .CK(clknet_leaf_181_clk),
    .Q(\g_row[0].g_col[1].mult.adder.b[9] ),
    .QN(_13437_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[0]$_DFF_PN0_  (.D(_00208_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.b[0] ),
    .QN(_00449_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[10]$_DFF_PN0_  (.D(_00209_),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_reduce0[0].adder.b[10] ),
    .QN(_00450_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[11]$_DFF_PN0_  (.D(_00210_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.b[11] ),
    .QN(_20359_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[12]$_DFF_PN0_  (.D(_00211_),
    .RN(net350),
    .CK(clknet_leaf_171_clk),
    .Q(\g_reduce0[0].adder.b[12] ),
    .QN(_20356_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[13]$_DFF_PN0_  (.D(_00212_),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_reduce0[0].adder.b[13] ),
    .QN(_20353_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[14]$_DFF_PN0_  (.D(_00213_),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_reduce0[0].adder.b[14] ),
    .QN(_20398_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[15]$_DFF_PN0_  (.D(\g_row[0].g_col[1].mult.sign ),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_reduce0[0].adder.b[15] ),
    .QN(_13438_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[1]$_DFF_PN0_  (.D(_00214_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[1] ),
    .QN(_20386_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[2]$_DFF_PN0_  (.D(_00215_),
    .RN(net276),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[2] ),
    .QN(_20383_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[3]$_DFF_PN0_  (.D(_00216_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[3] ),
    .QN(_20380_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[4]$_DFF_PN0_  (.D(_00217_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[4] ),
    .QN(_20377_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[5]$_DFF_PN0_  (.D(_00218_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[5] ),
    .QN(_20374_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[6]$_DFF_PN0_  (.D(_00219_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[6] ),
    .QN(_20371_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[7]$_DFF_PN0_  (.D(_00220_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.b[7] ),
    .QN(_20368_));
 DFFR_X2 \g_row[0].g_col[1].mult.x[8]$_DFF_PN0_  (.D(_00221_),
    .RN(net276),
    .CK(clknet_leaf_173_clk),
    .Q(\g_reduce0[0].adder.b[8] ),
    .QN(_20365_));
 DFFR_X1 \g_row[0].g_col[1].mult.x[9]$_DFF_PN0_  (.D(_00222_),
    .RN(net350),
    .CK(clknet_leaf_172_clk),
    .Q(\g_reduce0[0].adder.b[9] ),
    .QN(_20362_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.expa[0]$_DFF_PN0_  (.D(net173),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14255_));
 DFFR_X2 \g_row[0].g_col[2].mult.stage1.expa[1]$_DFF_PN0_  (.D(net174),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14260_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.expa[2]$_DFF_PN0_  (.D(net175),
    .RN(net346),
    .CK(clknet_leaf_111_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13439_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.expa[3]$_DFF_PN0_  (.D(net176),
    .RN(net346),
    .CK(clknet_leaf_111_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13440_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.expa[4]$_DFF_PN0_  (.D(net177),
    .RN(net346),
    .CK(clknet_leaf_111_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13441_));
 DFFR_X2 \g_row[0].g_col[2].mult.stage1.expb[0]$_DFF_PN0_  (.D(net256),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[0].fa.b ),
    .QN(_14254_));
 DFFR_X2 \g_row[0].g_col[2].mult.stage1.expb[1]$_DFF_PN0_  (.D(net257),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[1].fa.b ),
    .QN(_14259_));
 DFFR_X2 \g_row[0].g_col[2].mult.stage1.expb[2]$_DFF_PN0_  (.D(net258),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[2].fa.b ),
    .QN(_13442_));
 DFFR_X2 \g_row[0].g_col[2].mult.stage1.expb[3]$_DFF_PN0_  (.D(net259),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[3].fa.b ),
    .QN(_13443_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.expb[4]$_DFF_PN0_  (.D(net260),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[0].g_col[2].mult.expAdder.g_intermediate[4].fa.b ),
    .QN(_13444_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.sign$_DFF_PN0_  (.D(_00239_),
    .RN(net349),
    .CK(clknet_leaf_109_clk),
    .Q(\g_row[0].g_col[2].mult.sign ),
    .QN(_13445_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[0] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[0] ),
    .QN(_13446_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[10] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[10] ),
    .QN(_13447_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[11] ),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[11] ),
    .QN(_13448_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[12] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[12] ),
    .QN(_13449_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[13] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[13] ),
    .QN(_13450_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[14] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[14] ),
    .QN(_13451_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[15] ),
    .RN(net346),
    .CK(clknet_leaf_84_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[15] ),
    .QN(_13452_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[16] ),
    .RN(net346),
    .CK(clknet_leaf_84_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[16] ),
    .QN(_13453_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[17] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[17] ),
    .QN(_13454_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[18] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[18] ),
    .QN(_13455_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[19] ),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[19] ),
    .QN(_13456_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[1] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[1] ),
    .QN(_13457_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[2] ),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[2] ),
    .QN(_14249_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[3] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[3] ),
    .QN(_13458_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[4] ),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[4] ),
    .QN(_13459_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[5] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[5] ),
    .QN(_13460_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[6] ),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[6] ),
    .QN(_13461_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[7] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[7] ),
    .QN(_13462_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[8] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[8] ),
    .QN(_13463_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t1[9] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.a[9] ),
    .QN(_13464_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[10] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[10] ),
    .QN(_13465_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[11] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[11] ),
    .QN(_13466_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[12] ),
    .RN(net346),
    .CK(clknet_leaf_84_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[12] ),
    .QN(_13467_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[13] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[13] ),
    .QN(_13468_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[14] ),
    .RN(net346),
    .CK(clknet_leaf_84_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[14] ),
    .QN(_13469_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[15] ),
    .RN(net346),
    .CK(clknet_leaf_84_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[15] ),
    .QN(_13470_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[16] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[16] ),
    .QN(_13471_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[17] ),
    .RN(net346),
    .CK(clknet_leaf_83_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[17] ),
    .QN(_13472_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[18] ),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[18] ),
    .QN(_13473_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[19] ),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[19] ),
    .QN(_13474_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[1] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[1] ),
    .QN(_13475_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[20] ),
    .RN(net346),
    .CK(clknet_leaf_75_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[20] ),
    .QN(_13476_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[2] ),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[2] ),
    .QN(_14250_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[3] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[3] ),
    .QN(_13477_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[4] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[4] ),
    .QN(_13478_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[5] ),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[5] ),
    .QN(_13479_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[6] ),
    .RN(net346),
    .CK(clknet_leaf_80_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[6] ),
    .QN(_13480_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[7] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[7] ),
    .QN(_13481_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[8] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[8] ),
    .QN(_13482_));
 DFFR_X1 \g_row[0].g_col[2].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.stage1.dadda.t2[9] ),
    .RN(net346),
    .CK(clknet_leaf_81_clk),
    .Q(\g_row[0].g_col[2].mult.adder.b[9] ),
    .QN(_13483_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[0]$_DFF_PN0_  (.D(_00224_),
    .RN(net349),
    .CK(clknet_leaf_117_clk),
    .Q(\g_reduce0[2].adder.a[0] ),
    .QN(_21445_));
 DFFR_X2 \g_row[0].g_col[2].mult.x[10]$_DFF_PN0_  (.D(_00225_),
    .RN(net349),
    .CK(clknet_leaf_117_clk),
    .Q(\g_reduce0[2].adder.a[10] ),
    .QN(_21448_));
 DFFR_X2 \g_row[0].g_col[2].mult.x[11]$_DFF_PN0_  (.D(_00226_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.a[11] ),
    .QN(_00509_));
 DFFR_X2 \g_row[0].g_col[2].mult.x[12]$_DFF_PN0_  (.D(_00227_),
    .RN(net349),
    .CK(clknet_leaf_113_clk),
    .Q(\g_reduce0[2].adder.a[12] ),
    .QN(_00514_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[13]$_DFF_PN0_  (.D(_00228_),
    .RN(net349),
    .CK(clknet_leaf_113_clk),
    .Q(\g_reduce0[2].adder.a[13] ),
    .QN(_00517_));
 DFFR_X2 \g_row[0].g_col[2].mult.x[14]$_DFF_PN0_  (.D(_00229_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.a[14] ),
    .QN(_13484_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[15]$_DFF_PN0_  (.D(\g_row[0].g_col[2].mult.sign ),
    .RN(net348),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[2].adder.a[15] ),
    .QN(_13485_));
 DFFR_X2 \g_row[0].g_col[2].mult.x[1]$_DFF_PN0_  (.D(_00230_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[1] ),
    .QN(_00504_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[2]$_DFF_PN0_  (.D(_00231_),
    .RN(net349),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[2].adder.a[2] ),
    .QN(_00508_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[3]$_DFF_PN0_  (.D(_00232_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[3] ),
    .QN(_00507_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[4]$_DFF_PN0_  (.D(_00233_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[4] ),
    .QN(_00511_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[5]$_DFF_PN0_  (.D(_00234_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[5] ),
    .QN(_00510_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[6]$_DFF_PN0_  (.D(_00235_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[6] ),
    .QN(_00513_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[7]$_DFF_PN0_  (.D(_00236_),
    .RN(net349),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[2].adder.a[7] ),
    .QN(_00512_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[8]$_DFF_PN0_  (.D(_00237_),
    .RN(net349),
    .CK(clknet_leaf_115_clk),
    .Q(\g_reduce0[2].adder.a[8] ),
    .QN(_00516_));
 DFFR_X1 \g_row[0].g_col[2].mult.x[9]$_DFF_PN0_  (.D(_00238_),
    .RN(net349),
    .CK(clknet_leaf_116_clk),
    .Q(\g_reduce0[2].adder.a[9] ),
    .QN(_00515_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.expa[0]$_DFF_PN0_  (.D(net188),
    .RN(net349),
    .CK(clknet_leaf_107_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14274_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expa[1]$_DFF_PN0_  (.D(net189),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14279_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expa[2]$_DFF_PN0_  (.D(net191),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13486_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expa[3]$_DFF_PN0_  (.D(net192),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13487_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expa[4]$_DFF_PN0_  (.D(net193),
    .RN(net346),
    .CK(clknet_leaf_98_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13488_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expb[0]$_DFF_PN0_  (.D(net268),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[0].fa.b ),
    .QN(_14273_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expb[1]$_DFF_PN0_  (.D(net269),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[1].fa.b ),
    .QN(_14278_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expb[2]$_DFF_PN0_  (.D(net271),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[2].fa.b ),
    .QN(_13489_));
 DFFR_X2 \g_row[0].g_col[3].mult.stage1.expb[3]$_DFF_PN0_  (.D(net272),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[3].fa.b ),
    .QN(_13490_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.expb[4]$_DFF_PN0_  (.D(net273),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[0].g_col[3].mult.expAdder.g_intermediate[4].fa.b ),
    .QN(_13491_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.sign$_DFF_PN0_  (.D(_00255_),
    .RN(net349),
    .CK(clknet_leaf_107_clk),
    .Q(\g_row[0].g_col[3].mult.sign ),
    .QN(_13492_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[0] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[0] ),
    .QN(_13493_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[10] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[10] ),
    .QN(_13494_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[11] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[11] ),
    .QN(_13495_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[12] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[12] ),
    .QN(_13496_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[13] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[13] ),
    .QN(_13497_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[14] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[14] ),
    .QN(_13498_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[15] ),
    .RN(net350),
    .CK(clknet_leaf_157_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[15] ),
    .QN(_13499_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[16] ),
    .RN(net350),
    .CK(clknet_leaf_157_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[16] ),
    .QN(_13500_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[17] ),
    .RN(net350),
    .CK(clknet_leaf_157_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[17] ),
    .QN(_13501_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[18] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[18] ),
    .QN(_13502_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[19] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[19] ),
    .QN(_13503_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[1] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[1] ),
    .QN(_13504_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[2] ),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[2] ),
    .QN(_14268_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[3] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[3] ),
    .QN(_13505_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[4] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[4] ),
    .QN(_13506_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[5] ),
    .RN(net350),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[5] ),
    .QN(_13507_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[6] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[6] ),
    .QN(_13508_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[7] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[7] ),
    .QN(_13509_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[8] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[8] ),
    .QN(_13510_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t1[9] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.a[9] ),
    .QN(_13511_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[10] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[10] ),
    .QN(_13512_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[11] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[11] ),
    .QN(_13513_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[12] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[12] ),
    .QN(_13514_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[13] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[13] ),
    .QN(_13515_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[14] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[14] ),
    .QN(_13516_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[15] ),
    .RN(net350),
    .CK(clknet_leaf_157_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[15] ),
    .QN(_13517_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[16] ),
    .RN(net350),
    .CK(clknet_leaf_156_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[16] ),
    .QN(_13518_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[17] ),
    .RN(net350),
    .CK(clknet_leaf_157_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[17] ),
    .QN(_13519_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[18] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[18] ),
    .QN(_13520_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[19] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[19] ),
    .QN(_13521_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[1] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[1] ),
    .QN(_13522_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[20] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[20] ),
    .QN(_13523_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[2] ),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[2] ),
    .QN(_14269_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[3] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[3] ),
    .QN(_13524_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[4] ),
    .RN(net349),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[4] ),
    .QN(_13525_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[5] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[5] ),
    .QN(_13526_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[6] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[6] ),
    .QN(_13527_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[7] ),
    .RN(net350),
    .CK(clknet_leaf_154_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[7] ),
    .QN(_13528_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[8] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[8] ),
    .QN(_13529_));
 DFFR_X1 \g_row[0].g_col[3].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.stage1.dadda.t2[9] ),
    .RN(net350),
    .CK(clknet_leaf_155_clk),
    .Q(\g_row[0].g_col[3].mult.adder.b[9] ),
    .QN(_13530_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[0]$_DFF_PN0_  (.D(_00240_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[0] ),
    .QN(_00505_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[10]$_DFF_PN0_  (.D(_00241_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.b[10] ),
    .QN(_00506_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[11]$_DFF_PN0_  (.D(_00242_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.b[11] ),
    .QN(_21415_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[12]$_DFF_PN0_  (.D(_00243_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.b[12] ),
    .QN(_21412_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[13]$_DFF_PN0_  (.D(_00244_),
    .RN(net349),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[2].adder.b[13] ),
    .QN(_21409_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[14]$_DFF_PN0_  (.D(_00245_),
    .RN(net349),
    .CK(clknet_leaf_113_clk),
    .Q(\g_reduce0[2].adder.b[14] ),
    .QN(_21454_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[15]$_DFF_PN0_  (.D(\g_row[0].g_col[3].mult.sign ),
    .RN(net348),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[2].adder.b[15] ),
    .QN(_13531_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[1]$_DFF_PN0_  (.D(_00246_),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_reduce0[2].adder.b[1] ),
    .QN(_21442_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[2]$_DFF_PN0_  (.D(_00247_),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_reduce0[2].adder.b[2] ),
    .QN(_21439_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[3]$_DFF_PN0_  (.D(_00248_),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_reduce0[2].adder.b[3] ),
    .QN(_21436_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[4]$_DFF_PN0_  (.D(_00249_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[4] ),
    .QN(_21433_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[5]$_DFF_PN0_  (.D(_00250_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[5] ),
    .QN(_21430_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[6]$_DFF_PN0_  (.D(_00251_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[6] ),
    .QN(_21427_));
 DFFR_X2 \g_row[0].g_col[3].mult.x[7]$_DFF_PN0_  (.D(_00252_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[7] ),
    .QN(_21424_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[8]$_DFF_PN0_  (.D(_00253_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[8] ),
    .QN(_21421_));
 DFFR_X1 \g_row[0].g_col[3].mult.x[9]$_DFF_PN0_  (.D(_00254_),
    .RN(net349),
    .CK(clknet_leaf_158_clk),
    .Q(\g_reduce0[2].adder.b[9] ),
    .QN(_21418_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.expa[0]$_DFF_PN0_  (.D(net205),
    .RN(net347),
    .CK(clknet_leaf_27_clk),
    .Q(\g_row[1].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14292_));
 DFFR_X2 \g_row[1].g_col[0].mult.stage1.expa[1]$_DFF_PN0_  (.D(net206),
    .RN(net347),
    .CK(clknet_leaf_27_clk),
    .Q(\g_row[1].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14296_));
 DFFR_X2 \g_row[1].g_col[0].mult.stage1.expa[2]$_DFF_PN0_  (.D(net207),
    .RN(net351),
    .CK(clknet_leaf_39_clk),
    .Q(\g_row[1].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13532_));
 DFFR_X2 \g_row[1].g_col[0].mult.stage1.expa[3]$_DFF_PN0_  (.D(net208),
    .RN(net351),
    .CK(clknet_leaf_38_clk),
    .Q(\g_row[1].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13533_));
 DFFR_X2 \g_row[1].g_col[0].mult.stage1.expa[4]$_DFF_PN0_  (.D(net209),
    .RN(net351),
    .CK(clknet_leaf_38_clk),
    .Q(\g_row[1].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13534_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.sign$_DFF_PN0_  (.D(_00271_),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_row[1].g_col[0].mult.sign ),
    .QN(_13535_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[0] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[0] ),
    .QN(_13536_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[10] ),
    .RN(net345),
    .CK(clknet_leaf_51_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[10] ),
    .QN(_13537_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[11] ),
    .RN(net345),
    .CK(clknet_leaf_51_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[11] ),
    .QN(_13538_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[12] ),
    .RN(net345),
    .CK(clknet_leaf_51_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[12] ),
    .QN(_13539_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[13] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[13] ),
    .QN(_13540_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[14] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[14] ),
    .QN(_13541_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[15] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[15] ),
    .QN(_13542_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[16] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[16] ),
    .QN(_13543_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[17] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[17] ),
    .QN(_13544_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[18] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[18] ),
    .QN(_13545_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[19] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[19] ),
    .QN(_13546_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[1] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[1] ),
    .QN(_13547_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[2] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[2] ),
    .QN(_14287_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[3] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[3] ),
    .QN(_13548_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[4] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[4] ),
    .QN(_13549_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[5] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[5] ),
    .QN(_13550_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[6] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[6] ),
    .QN(_13551_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[7] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[7] ),
    .QN(_13552_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[8] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[8] ),
    .QN(_13553_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t1[9] ),
    .RN(net345),
    .CK(clknet_leaf_51_clk),
    .Q(\g_row[1].g_col[0].mult.adder.a[9] ),
    .QN(_13554_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[10] ),
    .RN(net345),
    .CK(clknet_leaf_51_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[10] ),
    .QN(_13555_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[11] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[11] ),
    .QN(_13556_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[12] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[12] ),
    .QN(_13557_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[13] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[13] ),
    .QN(_13558_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[14] ),
    .RN(net345),
    .CK(clknet_leaf_50_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[14] ),
    .QN(_13559_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[15] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[15] ),
    .QN(_13560_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[16] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[16] ),
    .QN(_13561_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[17] ),
    .RN(net345),
    .CK(clknet_leaf_49_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[17] ),
    .QN(_13562_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[18] ),
    .RN(net345),
    .CK(clknet_leaf_49_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[18] ),
    .QN(_13563_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[19] ),
    .RN(net345),
    .CK(clknet_leaf_48_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[19] ),
    .QN(_13564_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[1] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[1] ),
    .QN(_13565_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[20] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[20] ),
    .QN(_13566_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[2] ),
    .RN(net345),
    .CK(clknet_leaf_54_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[2] ),
    .QN(_14288_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[3] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[3] ),
    .QN(_13567_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[4] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[4] ),
    .QN(_13568_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[5] ),
    .RN(net345),
    .CK(clknet_leaf_53_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[5] ),
    .QN(_13569_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[6] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[6] ),
    .QN(_13570_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[7] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[7] ),
    .QN(_13571_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[8] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[8] ),
    .QN(_13572_));
 DFFR_X1 \g_row[1].g_col[0].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.stage1.dadda.t2[9] ),
    .RN(net345),
    .CK(clknet_leaf_52_clk),
    .Q(\g_row[1].g_col[0].mult.adder.b[9] ),
    .QN(_13573_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[0]$_DFF_PN0_  (.D(_00256_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.a[0] ),
    .QN(_00520_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[10]$_DFF_PN0_  (.D(_00257_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.a[10] ),
    .QN(_13574_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[11]$_DFF_PN0_  (.D(_00258_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.a[11] ),
    .QN(_21562_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[12]$_DFF_PN0_  (.D(_00259_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.a[12] ),
    .QN(_21559_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[13]$_DFF_PN0_  (.D(_00260_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.a[13] ),
    .QN(_21556_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[14]$_DFF_PN0_  (.D(_00261_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.a[14] ),
    .QN(_21598_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[15]$_DFF_PN0_  (.D(\g_row[1].g_col[0].mult.sign ),
    .RN(net347),
    .CK(clknet_leaf_160_clk),
    .Q(\g_reduce0[4].adder.a[15] ),
    .QN(_13575_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[1]$_DFF_PN0_  (.D(_00262_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.a[1] ),
    .QN(_21592_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[2]$_DFF_PN0_  (.D(_00263_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.a[2] ),
    .QN(_21589_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[3]$_DFF_PN0_  (.D(_00264_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.a[3] ),
    .QN(_21586_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[4]$_DFF_PN0_  (.D(_00265_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.a[4] ),
    .QN(_21583_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[5]$_DFF_PN0_  (.D(_00266_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[4].adder.a[5] ),
    .QN(_21580_));
 DFFR_X1 \g_row[1].g_col[0].mult.x[6]$_DFF_PN0_  (.D(_00267_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.a[6] ),
    .QN(_21577_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[7]$_DFF_PN0_  (.D(_00268_),
    .RN(net347),
    .CK(clknet_leaf_24_clk),
    .Q(\g_reduce0[4].adder.a[7] ),
    .QN(_21574_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[8]$_DFF_PN0_  (.D(_00269_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.a[8] ),
    .QN(_21571_));
 DFFR_X2 \g_row[1].g_col[0].mult.x[9]$_DFF_PN0_  (.D(_00270_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.a[9] ),
    .QN(_21568_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.expa[0]$_DFF_PN0_  (.D(net222),
    .RN(net276),
    .CK(clknet_leaf_20_clk),
    .Q(\g_row[1].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14309_));
 DFFR_X2 \g_row[1].g_col[1].mult.stage1.expa[1]$_DFF_PN0_  (.D(net223),
    .RN(net276),
    .CK(clknet_leaf_20_clk),
    .Q(\g_row[1].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14313_));
 DFFR_X2 \g_row[1].g_col[1].mult.stage1.expa[2]$_DFF_PN0_  (.D(net224),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[1].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13576_));
 DFFR_X2 \g_row[1].g_col[1].mult.stage1.expa[3]$_DFF_PN0_  (.D(net225),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_row[1].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13577_));
 DFFR_X2 \g_row[1].g_col[1].mult.stage1.expa[4]$_DFF_PN0_  (.D(net226),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[1].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13578_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.sign$_DFF_PN0_  (.D(_00287_),
    .RN(net350),
    .CK(clknet_leaf_166_clk),
    .Q(\g_row[1].g_col[1].mult.sign ),
    .QN(_13579_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[0] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[0] ),
    .QN(_13580_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[10] ),
    .RN(net276),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[10] ),
    .QN(_13581_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[11] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[11] ),
    .QN(_13582_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[12] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[12] ),
    .QN(_13583_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[13] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[13] ),
    .QN(_13584_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[14] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[14] ),
    .QN(_13585_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[15] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[15] ),
    .QN(_13586_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[16] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[16] ),
    .QN(_13587_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[17] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[17] ),
    .QN(_13588_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[18] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[18] ),
    .QN(_13589_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[19] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[19] ),
    .QN(_13590_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[1] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[1] ),
    .QN(_13591_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[2] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[2] ),
    .QN(_14304_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[3] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[3] ),
    .QN(_13592_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[4] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[4] ),
    .QN(_13593_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[5] ),
    .RN(net276),
    .CK(clknet_leaf_4_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[5] ),
    .QN(_13594_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[6] ),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[6] ),
    .QN(_13595_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[7] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[7] ),
    .QN(_13596_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[8] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[8] ),
    .QN(_13597_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t1[9] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.a[9] ),
    .QN(_13598_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[10] ),
    .RN(net276),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[10] ),
    .QN(_13599_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[11] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[11] ),
    .QN(_13600_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[12] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[12] ),
    .QN(_13601_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[13] ),
    .RN(net347),
    .CK(clknet_leaf_15_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[13] ),
    .QN(_13602_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[14] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[14] ),
    .QN(_13603_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[15] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[15] ),
    .QN(_13604_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[16] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[16] ),
    .QN(_13605_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[17] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[17] ),
    .QN(_13606_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[18] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[18] ),
    .QN(_13607_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[19] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[19] ),
    .QN(_13608_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[1] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[1] ),
    .QN(_13609_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[20] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[20] ),
    .QN(_13610_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[2] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[2] ),
    .QN(_14305_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[3] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[3] ),
    .QN(_13611_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[4] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[4] ),
    .QN(_13612_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[5] ),
    .RN(net276),
    .CK(clknet_leaf_17_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[5] ),
    .QN(_13613_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[6] ),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[6] ),
    .QN(_13614_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[7] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[7] ),
    .QN(_13615_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[8] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[8] ),
    .QN(_13616_));
 DFFR_X1 \g_row[1].g_col[1].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.stage1.dadda.t2[9] ),
    .RN(net276),
    .CK(clknet_leaf_16_clk),
    .Q(\g_row[1].g_col[1].mult.adder.b[9] ),
    .QN(_13617_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[0]$_DFF_PN0_  (.D(_00272_),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_reduce0[4].adder.b[0] ),
    .QN(_00519_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[10]$_DFF_PN0_  (.D(_00273_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.b[10] ),
    .QN(_21565_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[11]$_DFF_PN0_  (.D(_00274_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.b[11] ),
    .QN(_00523_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[12]$_DFF_PN0_  (.D(_00275_),
    .RN(net347),
    .CK(clknet_leaf_25_clk),
    .Q(\g_reduce0[4].adder.b[12] ),
    .QN(_00528_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[13]$_DFF_PN0_  (.D(_00276_),
    .RN(net347),
    .CK(clknet_leaf_23_clk),
    .Q(\g_reduce0[4].adder.b[13] ),
    .QN(_00531_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[14]$_DFF_PN0_  (.D(_00277_),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_reduce0[4].adder.b[14] ),
    .QN(_13618_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[15]$_DFF_PN0_  (.D(\g_row[1].g_col[1].mult.sign ),
    .RN(net276),
    .CK(clknet_leaf_164_clk),
    .Q(\g_reduce0[4].adder.b[15] ),
    .QN(_13619_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[1]$_DFF_PN0_  (.D(_00278_),
    .RN(net347),
    .CK(clknet_leaf_26_clk),
    .Q(\g_reduce0[4].adder.b[1] ),
    .QN(_00518_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[2]$_DFF_PN0_  (.D(_00279_),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_reduce0[4].adder.b[2] ),
    .QN(_00522_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[3]$_DFF_PN0_  (.D(_00280_),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_reduce0[4].adder.b[3] ),
    .QN(_00521_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[4]$_DFF_PN0_  (.D(_00281_),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_reduce0[4].adder.b[4] ),
    .QN(_00525_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[5]$_DFF_PN0_  (.D(_00282_),
    .RN(net347),
    .CK(clknet_leaf_22_clk),
    .Q(\g_reduce0[4].adder.b[5] ),
    .QN(_00524_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[6]$_DFF_PN0_  (.D(_00283_),
    .RN(net347),
    .CK(clknet_leaf_22_clk),
    .Q(\g_reduce0[4].adder.b[6] ),
    .QN(_00527_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[7]$_DFF_PN0_  (.D(_00284_),
    .RN(net347),
    .CK(clknet_leaf_22_clk),
    .Q(\g_reduce0[4].adder.b[7] ),
    .QN(_00526_));
 DFFR_X2 \g_row[1].g_col[1].mult.x[8]$_DFF_PN0_  (.D(_00285_),
    .RN(net347),
    .CK(clknet_leaf_22_clk),
    .Q(\g_reduce0[4].adder.b[8] ),
    .QN(_00530_));
 DFFR_X1 \g_row[1].g_col[1].mult.x[9]$_DFF_PN0_  (.D(_00286_),
    .RN(net347),
    .CK(clknet_leaf_22_clk),
    .Q(\g_reduce0[4].adder.b[9] ),
    .QN(_00529_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.expa[0]$_DFF_PN0_  (.D(net6),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_row[1].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14326_));
 DFFR_X2 \g_row[1].g_col[2].mult.stage1.expa[1]$_DFF_PN0_  (.D(net7),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_row[1].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14331_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.expa[2]$_DFF_PN0_  (.D(net8),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_row[1].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13620_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.expa[3]$_DFF_PN0_  (.D(net9),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[1].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13621_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.expa[4]$_DFF_PN0_  (.D(net11),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_row[1].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13622_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.sign$_DFF_PN0_  (.D(_00303_),
    .RN(net348),
    .CK(clknet_leaf_105_clk),
    .Q(\g_row[1].g_col[2].mult.sign ),
    .QN(_13623_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[0] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[0] ),
    .QN(_13624_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[10] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[10] ),
    .QN(_13625_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[11] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[11] ),
    .QN(_13626_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[12] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[12] ),
    .QN(_13627_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[13] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[13] ),
    .QN(_13628_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[14] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[14] ),
    .QN(_13629_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[15] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[15] ),
    .QN(_13630_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[16] ),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[16] ),
    .QN(_13631_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[17] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[17] ),
    .QN(_13632_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[18] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[18] ),
    .QN(_13633_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[19] ),
    .RN(net345),
    .CK(clknet_leaf_85_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[19] ),
    .QN(_13634_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[1] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[1] ),
    .QN(_13635_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[2] ),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[2] ),
    .QN(_14321_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[3] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[3] ),
    .QN(_13636_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[4] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[4] ),
    .QN(_13637_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[5] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[5] ),
    .QN(_13638_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[6] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[6] ),
    .QN(_13639_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[7] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[7] ),
    .QN(_13640_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[8] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[8] ),
    .QN(_13641_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t1[9] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.a[9] ),
    .QN(_13642_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[10] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[10] ),
    .QN(_13643_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[11] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[11] ),
    .QN(_13644_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[12] ),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[12] ),
    .QN(_13645_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[13] ),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[13] ),
    .QN(_13646_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[14] ),
    .RN(net346),
    .CK(clknet_leaf_87_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[14] ),
    .QN(_13647_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[15] ),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[15] ),
    .QN(_13648_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[16] ),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[16] ),
    .QN(_13649_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[17] ),
    .RN(net346),
    .CK(clknet_leaf_88_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[17] ),
    .QN(_13650_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[18] ),
    .RN(net345),
    .CK(clknet_leaf_85_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[18] ),
    .QN(_13651_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[19] ),
    .RN(net345),
    .CK(clknet_leaf_85_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[19] ),
    .QN(_13652_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[1] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[1] ),
    .QN(_13653_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[20] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[20] ),
    .QN(_13654_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[2] ),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[2] ),
    .QN(_14322_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[3] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[3] ),
    .QN(_13655_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[4] ),
    .RN(net346),
    .CK(clknet_leaf_91_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[4] ),
    .QN(_13656_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[5] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[5] ),
    .QN(_13657_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[6] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[6] ),
    .QN(_13658_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[7] ),
    .RN(net346),
    .CK(clknet_leaf_90_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[7] ),
    .QN(_13659_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[8] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[8] ),
    .QN(_13660_));
 DFFR_X1 \g_row[1].g_col[2].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.stage1.dadda.t2[9] ),
    .RN(net346),
    .CK(clknet_leaf_86_clk),
    .Q(\g_row[1].g_col[2].mult.adder.b[9] ),
    .QN(_13661_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[0]$_DFF_PN0_  (.D(_00288_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.a[0] ),
    .QN(_21736_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[10]$_DFF_PN0_  (.D(_00289_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.a[10] ),
    .QN(_21739_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[11]$_DFF_PN0_  (.D(_00290_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.a[11] ),
    .QN(_00537_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[12]$_DFF_PN0_  (.D(_00291_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.a[12] ),
    .QN(_00542_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[13]$_DFF_PN0_  (.D(_00292_),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_reduce0[6].adder.a[13] ),
    .QN(_00545_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[14]$_DFF_PN0_  (.D(_00293_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.a[14] ),
    .QN(_13662_));
 DFFR_X2 \g_row[1].g_col[2].mult.x[15]$_DFF_PN0_  (.D(\g_row[1].g_col[2].mult.sign ),
    .RN(net346),
    .CK(clknet_leaf_101_clk),
    .Q(\g_reduce0[6].adder.a[15] ),
    .QN(_13663_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[1]$_DFF_PN0_  (.D(_00294_),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_reduce0[6].adder.a[1] ),
    .QN(_00532_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[2]$_DFF_PN0_  (.D(_00295_),
    .RN(net346),
    .CK(clknet_leaf_92_clk),
    .Q(\g_reduce0[6].adder.a[2] ),
    .QN(_00536_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[3]$_DFF_PN0_  (.D(_00296_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.a[3] ),
    .QN(_00535_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[4]$_DFF_PN0_  (.D(_00297_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.a[4] ),
    .QN(_00539_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[5]$_DFF_PN0_  (.D(_00298_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.a[5] ),
    .QN(_00538_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[6]$_DFF_PN0_  (.D(_00299_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.a[6] ),
    .QN(_00541_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[7]$_DFF_PN0_  (.D(_00300_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.a[7] ),
    .QN(_00540_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[8]$_DFF_PN0_  (.D(_00301_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.a[8] ),
    .QN(_00544_));
 DFFR_X1 \g_row[1].g_col[2].mult.x[9]$_DFF_PN0_  (.D(_00302_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.a[9] ),
    .QN(_00543_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.expa[0]$_DFF_PN0_  (.D(net22),
    .RN(net346),
    .CK(clknet_leaf_93_clk),
    .Q(\g_row[1].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14343_));
 DFFR_X2 \g_row[1].g_col[3].mult.stage1.expa[1]$_DFF_PN0_  (.D(net23),
    .RN(net346),
    .CK(clknet_leaf_93_clk),
    .Q(\g_row[1].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14348_));
 DFFR_X2 \g_row[1].g_col[3].mult.stage1.expa[2]$_DFF_PN0_  (.D(net24),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[1].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13664_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.expa[3]$_DFF_PN0_  (.D(net25),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[1].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13665_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.expa[4]$_DFF_PN0_  (.D(net26),
    .RN(net346),
    .CK(clknet_leaf_89_clk),
    .Q(\g_row[1].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13666_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.sign$_DFF_PN0_  (.D(_00319_),
    .RN(net348),
    .CK(clknet_leaf_105_clk),
    .Q(\g_row[1].g_col[3].mult.sign ),
    .QN(_13667_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[0] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[0] ),
    .QN(_13668_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[10] ),
    .RN(net349),
    .CK(clknet_leaf_149_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[10] ),
    .QN(_13669_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[11] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[11] ),
    .QN(_13670_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[12] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[12] ),
    .QN(_13671_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[13] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[13] ),
    .QN(_13672_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[14] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[14] ),
    .QN(_13673_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[15] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[15] ),
    .QN(_13674_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[16] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[16] ),
    .QN(_13675_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[17] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[17] ),
    .QN(_13676_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[18] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[18] ),
    .QN(_13677_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[19] ),
    .RN(net349),
    .CK(clknet_leaf_117_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[19] ),
    .QN(_13678_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[1] ),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[1] ),
    .QN(_13679_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[2] ),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[2] ),
    .QN(_14338_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[3] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[3] ),
    .QN(_13680_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[4] ),
    .RN(net348),
    .CK(clknet_leaf_139_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[4] ),
    .QN(_13681_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[5] ),
    .RN(net348),
    .CK(clknet_leaf_139_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[5] ),
    .QN(_13682_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[6] ),
    .RN(net348),
    .CK(clknet_leaf_128_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[6] ),
    .QN(_13683_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[7] ),
    .RN(net349),
    .CK(clknet_leaf_139_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[7] ),
    .QN(_13684_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[8] ),
    .RN(net349),
    .CK(clknet_leaf_139_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[8] ),
    .QN(_13685_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t1[9] ),
    .RN(net349),
    .CK(clknet_leaf_149_clk),
    .Q(\g_row[1].g_col[3].mult.adder.a[9] ),
    .QN(_13686_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[10] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[10] ),
    .QN(_13687_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[11] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[11] ),
    .QN(_13688_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[12] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[12] ),
    .QN(_13689_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[13] ),
    .RN(net349),
    .CK(clknet_leaf_151_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[13] ),
    .QN(_13690_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[14] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[14] ),
    .QN(_13691_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[15] ),
    .RN(net349),
    .CK(clknet_leaf_150_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[15] ),
    .QN(_13692_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[16] ),
    .RN(net349),
    .CK(clknet_leaf_118_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[16] ),
    .QN(_13693_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[17] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[17] ),
    .QN(_13694_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[18] ),
    .RN(net349),
    .CK(clknet_leaf_152_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[18] ),
    .QN(_13695_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[19] ),
    .RN(net349),
    .CK(clknet_leaf_117_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[19] ),
    .QN(_13696_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[1] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[1] ),
    .QN(_13697_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[20] ),
    .RN(net349),
    .CK(clknet_leaf_153_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[20] ),
    .QN(_13698_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[2] ),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[2] ),
    .QN(_14339_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[3] ),
    .RN(net348),
    .CK(clknet_leaf_138_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[3] ),
    .QN(_13699_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[4] ),
    .RN(net348),
    .CK(clknet_leaf_139_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[4] ),
    .QN(_13700_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[5] ),
    .RN(net348),
    .CK(clknet_leaf_128_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[5] ),
    .QN(_13701_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[6] ),
    .RN(net348),
    .CK(clknet_leaf_128_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[6] ),
    .QN(_13702_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[7] ),
    .RN(net349),
    .CK(clknet_leaf_128_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[7] ),
    .QN(_13703_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[8] ),
    .RN(net349),
    .CK(clknet_leaf_128_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[8] ),
    .QN(_13704_));
 DFFR_X1 \g_row[1].g_col[3].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.stage1.dadda.t2[9] ),
    .RN(net349),
    .CK(clknet_leaf_149_clk),
    .Q(\g_row[1].g_col[3].mult.adder.b[9] ),
    .QN(_13705_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[0]$_DFF_PN0_  (.D(_00304_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.b[0] ),
    .QN(_00533_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[10]$_DFF_PN0_  (.D(_00305_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.b[10] ),
    .QN(_00534_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[11]$_DFF_PN0_  (.D(_00306_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.b[11] ),
    .QN(_21706_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[12]$_DFF_PN0_  (.D(_00307_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.b[12] ),
    .QN(_21703_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[13]$_DFF_PN0_  (.D(_00308_),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_reduce0[6].adder.b[13] ),
    .QN(_21700_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[14]$_DFF_PN0_  (.D(_00309_),
    .RN(net346),
    .CK(clknet_leaf_96_clk),
    .Q(\g_reduce0[6].adder.b[14] ),
    .QN(_21745_));
 DFFR_X2 \g_row[1].g_col[3].mult.x[15]$_DFF_PN0_  (.D(\g_row[1].g_col[3].mult.sign ),
    .RN(net346),
    .CK(clknet_leaf_100_clk),
    .Q(\g_reduce0[6].adder.b[15] ),
    .QN(_13706_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[1]$_DFF_PN0_  (.D(_00310_),
    .RN(net346),
    .CK(clknet_leaf_93_clk),
    .Q(\g_reduce0[6].adder.b[1] ),
    .QN(_21733_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[2]$_DFF_PN0_  (.D(_00311_),
    .RN(net346),
    .CK(clknet_leaf_103_clk),
    .Q(\g_reduce0[6].adder.b[2] ),
    .QN(_21730_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[3]$_DFF_PN0_  (.D(_00312_),
    .RN(net346),
    .CK(clknet_leaf_102_clk),
    .Q(\g_reduce0[6].adder.b[3] ),
    .QN(_21727_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[4]$_DFF_PN0_  (.D(_00313_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.b[4] ),
    .QN(_21724_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[5]$_DFF_PN0_  (.D(_00314_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.b[5] ),
    .QN(_21721_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[6]$_DFF_PN0_  (.D(_00315_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.b[6] ),
    .QN(_21718_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[7]$_DFF_PN0_  (.D(_00316_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.b[7] ),
    .QN(_21715_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[8]$_DFF_PN0_  (.D(_00317_),
    .RN(net346),
    .CK(clknet_leaf_95_clk),
    .Q(\g_reduce0[6].adder.b[8] ),
    .QN(_21712_));
 DFFR_X1 \g_row[1].g_col[3].mult.x[9]$_DFF_PN0_  (.D(_00318_),
    .RN(net346),
    .CK(clknet_leaf_94_clk),
    .Q(\g_reduce0[6].adder.b[9] ),
    .QN(_21709_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.expa[0]$_DFF_PN0_  (.D(net37),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[2].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14360_));
 DFFR_X2 \g_row[2].g_col[0].mult.stage1.expa[1]$_DFF_PN0_  (.D(net38),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[2].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14364_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.expa[2]$_DFF_PN0_  (.D(net40),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[2].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13707_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.expa[3]$_DFF_PN0_  (.D(net41),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[2].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13708_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.expa[4]$_DFF_PN0_  (.D(net42),
    .RN(net351),
    .CK(clknet_leaf_34_clk),
    .Q(\g_row[2].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13709_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.sign$_DFF_PN0_  (.D(_00335_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_row[2].g_col[0].mult.sign ),
    .QN(_13710_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[0] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[0] ),
    .QN(_13711_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[10] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[10] ),
    .QN(_13712_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[11] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[11] ),
    .QN(_13713_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[12] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[12] ),
    .QN(_13714_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[13] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[13] ),
    .QN(_13715_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[14] ),
    .RN(net345),
    .CK(clknet_leaf_45_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[14] ),
    .QN(_13716_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[15] ),
    .RN(net345),
    .CK(clknet_leaf_45_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[15] ),
    .QN(_13717_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[16] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[16] ),
    .QN(_13718_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[17] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[17] ),
    .QN(_13719_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[18] ),
    .RN(net345),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[18] ),
    .QN(_13720_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[19] ),
    .RN(net345),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[19] ),
    .QN(_13721_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[1] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[1] ),
    .QN(_13722_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[2] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[2] ),
    .QN(_14355_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[3] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[3] ),
    .QN(_13723_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[4] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[4] ),
    .QN(_13724_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[5] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[5] ),
    .QN(_13725_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[6] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[6] ),
    .QN(_13726_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[7] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[7] ),
    .QN(_13727_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[8] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[8] ),
    .QN(_13728_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t1[9] ),
    .RN(net345),
    .CK(clknet_leaf_49_clk),
    .Q(\g_row[2].g_col[0].mult.adder.a[9] ),
    .QN(_13729_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[10] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[10] ),
    .QN(_13730_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[11] ),
    .RN(net345),
    .CK(clknet_leaf_49_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[11] ),
    .QN(_13731_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[12] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[12] ),
    .QN(_13732_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[13] ),
    .RN(net345),
    .CK(clknet_leaf_49_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[13] ),
    .QN(_13733_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[14] ),
    .RN(net345),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[14] ),
    .QN(_13734_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[15] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[15] ),
    .QN(_13735_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[16] ),
    .RN(net345),
    .CK(clknet_leaf_45_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[16] ),
    .QN(_13736_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[17] ),
    .RN(net345),
    .CK(clknet_leaf_42_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[17] ),
    .QN(_13737_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[18] ),
    .RN(net345),
    .CK(clknet_leaf_41_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[18] ),
    .QN(_13738_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[19] ),
    .RN(net345),
    .CK(clknet_leaf_45_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[19] ),
    .QN(_13739_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[1] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[1] ),
    .QN(_13740_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[20] ),
    .RN(net351),
    .CK(clknet_leaf_44_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[20] ),
    .QN(_13741_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[2] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[2] ),
    .QN(_14356_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[3] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[3] ),
    .QN(_13742_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[4] ),
    .RN(net345),
    .CK(clknet_leaf_55_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[4] ),
    .QN(_13743_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[5] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[5] ),
    .QN(_13744_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[6] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[6] ),
    .QN(_13745_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[7] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[7] ),
    .QN(_13746_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[8] ),
    .RN(net345),
    .CK(clknet_leaf_47_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[8] ),
    .QN(_13747_));
 DFFR_X1 \g_row[2].g_col[0].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.stage1.dadda.t2[9] ),
    .RN(net345),
    .CK(clknet_leaf_46_clk),
    .Q(\g_row[2].g_col[0].mult.adder.b[9] ),
    .QN(_13748_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[0]$_DFF_PN0_  (.D(_00320_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.a[0] ),
    .QN(_00548_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[10]$_DFF_PN0_  (.D(_00321_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.a[10] ),
    .QN(_13749_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[11]$_DFF_PN0_  (.D(_00322_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.a[11] ),
    .QN(_21853_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[12]$_DFF_PN0_  (.D(_00323_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.a[12] ),
    .QN(_21850_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[13]$_DFF_PN0_  (.D(_00324_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.a[13] ),
    .QN(_21847_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[14]$_DFF_PN0_  (.D(_00325_),
    .RN(net351),
    .CK(clknet_leaf_27_clk),
    .Q(\g_reduce0[8].adder.a[14] ),
    .QN(_21889_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[15]$_DFF_PN0_  (.D(\g_row[2].g_col[0].mult.sign ),
    .RN(net351),
    .CK(clknet_leaf_29_clk),
    .Q(\g_reduce0[8].adder.a[15] ),
    .QN(_13750_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[1]$_DFF_PN0_  (.D(_00326_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.a[1] ),
    .QN(_21883_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[2]$_DFF_PN0_  (.D(_00327_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.a[2] ),
    .QN(_21880_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[3]$_DFF_PN0_  (.D(_00328_),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_reduce0[8].adder.a[3] ),
    .QN(_21877_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[4]$_DFF_PN0_  (.D(_00329_),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_reduce0[8].adder.a[4] ),
    .QN(_21874_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[5]$_DFF_PN0_  (.D(_00330_),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_reduce0[8].adder.a[5] ),
    .QN(_21871_));
 DFFR_X1 \g_row[2].g_col[0].mult.x[6]$_DFF_PN0_  (.D(_00331_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.a[6] ),
    .QN(_21868_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[7]$_DFF_PN0_  (.D(_00332_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.a[7] ),
    .QN(_21865_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[8]$_DFF_PN0_  (.D(_00333_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.a[8] ),
    .QN(_21862_));
 DFFR_X2 \g_row[2].g_col[0].mult.x[9]$_DFF_PN0_  (.D(_00334_),
    .RN(net351),
    .CK(clknet_leaf_29_clk),
    .Q(\g_reduce0[8].adder.a[9] ),
    .QN(_21859_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.expa[0]$_DFF_PN0_  (.D(net54),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_row[2].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14377_));
 DFFR_X2 \g_row[2].g_col[1].mult.stage1.expa[1]$_DFF_PN0_  (.D(net55),
    .RN(net347),
    .CK(clknet_leaf_21_clk),
    .Q(\g_row[2].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14381_));
 DFFR_X2 \g_row[2].g_col[1].mult.stage1.expa[2]$_DFF_PN0_  (.D(net56),
    .RN(net350),
    .CK(clknet_leaf_179_clk),
    .Q(\g_row[2].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13751_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.expa[3]$_DFF_PN0_  (.D(net57),
    .RN(net347),
    .CK(clknet_leaf_27_clk),
    .Q(\g_row[2].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13752_));
 DFFR_X2 \g_row[2].g_col[1].mult.stage1.expa[4]$_DFF_PN0_  (.D(net58),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[2].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13753_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.sign$_DFF_PN0_  (.D(_00351_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_row[2].g_col[1].mult.sign ),
    .QN(_13754_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[0] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[0] ),
    .QN(_13755_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[10] ),
    .RN(net347),
    .CK(clknet_leaf_4_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[10] ),
    .QN(_13756_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[11] ),
    .RN(net347),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[11] ),
    .QN(_13757_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[12] ),
    .RN(net347),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[12] ),
    .QN(_13758_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[13] ),
    .RN(net351),
    .CK(clknet_leaf_4_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[13] ),
    .QN(_13759_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[14] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[14] ),
    .QN(_13760_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[15] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[15] ),
    .QN(_13761_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[16] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[16] ),
    .QN(_13762_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[17] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[17] ),
    .QN(_13763_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[18] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[18] ),
    .QN(_13764_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[19] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[19] ),
    .QN(_13765_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[1] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[1] ),
    .QN(_13766_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[2] ),
    .RN(net347),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[2] ),
    .QN(_14372_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[3] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[3] ),
    .QN(_13767_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[4] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[4] ),
    .QN(_13768_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[5] ),
    .RN(net347),
    .CK(clknet_leaf_10_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[5] ),
    .QN(_13769_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[6] ),
    .RN(net347),
    .CK(clknet_leaf_10_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[6] ),
    .QN(_13770_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[7] ),
    .RN(net347),
    .CK(clknet_leaf_10_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[7] ),
    .QN(_13771_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[8] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[8] ),
    .QN(_13772_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t1[9] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.a[9] ),
    .QN(_13773_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[10] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[10] ),
    .QN(_13774_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[11] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[11] ),
    .QN(_13775_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[12] ),
    .RN(net347),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[12] ),
    .QN(_13776_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[13] ),
    .RN(net351),
    .CK(clknet_leaf_4_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[13] ),
    .QN(_13777_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[14] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[14] ),
    .QN(_13778_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[15] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[15] ),
    .QN(_13779_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[16] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[16] ),
    .QN(_13780_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[17] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[17] ),
    .QN(_13781_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[18] ),
    .RN(net351),
    .CK(clknet_leaf_6_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[18] ),
    .QN(_13782_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[19] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[19] ),
    .QN(_13783_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[1] ),
    .RN(net347),
    .CK(clknet_leaf_13_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[1] ),
    .QN(_13784_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[20] ),
    .RN(net351),
    .CK(clknet_leaf_7_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[20] ),
    .QN(_13785_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[2] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[2] ),
    .QN(_14373_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[3] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[3] ),
    .QN(_13786_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[4] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[4] ),
    .QN(_13787_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[5] ),
    .RN(net347),
    .CK(clknet_leaf_14_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[5] ),
    .QN(_13788_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[6] ),
    .RN(net347),
    .CK(clknet_leaf_10_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[6] ),
    .QN(_13789_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[7] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[7] ),
    .QN(_13790_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[8] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[8] ),
    .QN(_13791_));
 DFFR_X1 \g_row[2].g_col[1].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.stage1.dadda.t2[9] ),
    .RN(net347),
    .CK(clknet_leaf_5_clk),
    .Q(\g_row[2].g_col[1].mult.adder.b[9] ),
    .QN(_13792_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[0]$_DFF_PN0_  (.D(_00336_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.b[0] ),
    .QN(_00547_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[10]$_DFF_PN0_  (.D(_00337_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.b[10] ),
    .QN(_21856_));
 DFFR_X2 \g_row[2].g_col[1].mult.x[11]$_DFF_PN0_  (.D(_00338_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.b[11] ),
    .QN(_00551_));
 DFFR_X2 \g_row[2].g_col[1].mult.x[12]$_DFF_PN0_  (.D(_00339_),
    .RN(net351),
    .CK(clknet_leaf_28_clk),
    .Q(\g_reduce0[8].adder.b[12] ),
    .QN(_00556_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[13]$_DFF_PN0_  (.D(_00340_),
    .RN(net351),
    .CK(clknet_leaf_29_clk),
    .Q(\g_reduce0[8].adder.b[13] ),
    .QN(_00559_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[14]$_DFF_PN0_  (.D(_00341_),
    .RN(net351),
    .CK(clknet_leaf_27_clk),
    .Q(\g_reduce0[8].adder.b[14] ),
    .QN(_13793_));
 DFFR_X2 \g_row[2].g_col[1].mult.x[15]$_DFF_PN0_  (.D(\g_row[2].g_col[1].mult.sign ),
    .RN(net351),
    .CK(clknet_leaf_27_clk),
    .Q(\g_reduce0[8].adder.b[15] ),
    .QN(_13794_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[1]$_DFF_PN0_  (.D(_00342_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.b[1] ),
    .QN(_00546_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[2]$_DFF_PN0_  (.D(_00343_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.b[2] ),
    .QN(_00550_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[3]$_DFF_PN0_  (.D(_00344_),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_reduce0[8].adder.b[3] ),
    .QN(_00549_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[4]$_DFF_PN0_  (.D(_00345_),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_reduce0[8].adder.b[4] ),
    .QN(_00553_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[5]$_DFF_PN0_  (.D(_00346_),
    .RN(net351),
    .CK(clknet_leaf_33_clk),
    .Q(\g_reduce0[8].adder.b[5] ),
    .QN(_00552_));
 DFFR_X2 \g_row[2].g_col[1].mult.x[6]$_DFF_PN0_  (.D(_00347_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.b[6] ),
    .QN(_00555_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[7]$_DFF_PN0_  (.D(_00348_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.b[7] ),
    .QN(_00554_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[8]$_DFF_PN0_  (.D(_00349_),
    .RN(net351),
    .CK(clknet_leaf_30_clk),
    .Q(\g_reduce0[8].adder.b[8] ),
    .QN(_00558_));
 DFFR_X1 \g_row[2].g_col[1].mult.x[9]$_DFF_PN0_  (.D(_00350_),
    .RN(net351),
    .CK(clknet_leaf_29_clk),
    .Q(\g_reduce0[8].adder.b[9] ),
    .QN(_00557_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.expa[0]$_DFF_PN0_  (.D(net70),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(\g_row[2].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14394_));
 DFFR_X2 \g_row[2].g_col[2].mult.stage1.expa[1]$_DFF_PN0_  (.D(net71),
    .RN(net346),
    .CK(clknet_leaf_77_clk),
    .Q(\g_row[2].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14399_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.expa[2]$_DFF_PN0_  (.D(net72),
    .RN(net346),
    .CK(clknet_leaf_82_clk),
    .Q(\g_row[2].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13795_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.expa[3]$_DFF_PN0_  (.D(net73),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[2].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13796_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.expa[4]$_DFF_PN0_  (.D(net74),
    .RN(net346),
    .CK(clknet_leaf_79_clk),
    .Q(\g_row[2].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13797_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.sign$_DFF_PN0_  (.D(_00367_),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[2].g_col[2].mult.sign ),
    .QN(_13798_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[0] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[0] ),
    .QN(_13799_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[10] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[10] ),
    .QN(_13800_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[11] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[11] ),
    .QN(_13801_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[12] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[12] ),
    .QN(_13802_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[13] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[13] ),
    .QN(_13803_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[14] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[14] ),
    .QN(_13804_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[15] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[15] ),
    .QN(_13805_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[16] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[16] ),
    .QN(_13806_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[17] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[17] ),
    .QN(_13807_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[18] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[18] ),
    .QN(_13808_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[19] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[19] ),
    .QN(_13809_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[1] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[1] ),
    .QN(_13810_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[2] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[2] ),
    .QN(_14389_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[3] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[3] ),
    .QN(_13811_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[4] ),
    .RN(net345),
    .CK(clknet_leaf_63_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[4] ),
    .QN(_13812_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[5] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[5] ),
    .QN(_13813_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[6] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[6] ),
    .QN(_13814_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[7] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[7] ),
    .QN(_13815_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[8] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[8] ),
    .QN(_13816_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t1[9] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.a[9] ),
    .QN(_13817_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[10] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[10] ),
    .QN(_13818_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[11] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[11] ),
    .QN(_13819_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[12] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[12] ),
    .QN(_13820_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[13] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[13] ),
    .QN(_13821_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[14] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[14] ),
    .QN(_13822_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[15] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[15] ),
    .QN(_13823_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[16] ),
    .RN(net345),
    .CK(clknet_leaf_58_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[16] ),
    .QN(_13824_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[17] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[17] ),
    .QN(_13825_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[18] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[18] ),
    .QN(_13826_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[19] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[19] ),
    .QN(_13827_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[1] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[1] ),
    .QN(_13828_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[20] ),
    .RN(net345),
    .CK(clknet_leaf_59_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[20] ),
    .QN(_13829_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[2] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[2] ),
    .QN(_14390_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[3] ),
    .RN(net345),
    .CK(clknet_leaf_62_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[3] ),
    .QN(_13830_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[4] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[4] ),
    .QN(_13831_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[5] ),
    .RN(net345),
    .CK(clknet_leaf_63_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[5] ),
    .QN(_13832_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[6] ),
    .RN(net345),
    .CK(clknet_leaf_63_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[6] ),
    .QN(_13833_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[7] ),
    .RN(net345),
    .CK(clknet_leaf_61_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[7] ),
    .QN(_13834_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[8] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[8] ),
    .QN(_13835_));
 DFFR_X1 \g_row[2].g_col[2].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.stage1.dadda.t2[9] ),
    .RN(net345),
    .CK(clknet_leaf_60_clk),
    .Q(\g_row[2].g_col[2].mult.adder.b[9] ),
    .QN(_13836_));
 DFFR_X1 \g_row[2].g_col[2].mult.x[0]$_DFF_PN0_  (.D(_00352_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.a[0] ),
    .QN(_00464_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[10]$_DFF_PN0_  (.D(_00353_),
    .RN(net346),
    .CK(clknet_leaf_76_clk),
    .Q(\g_reduce0[10].adder.a[10] ),
    .QN(_13837_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[11]$_DFF_PN0_  (.D(_00354_),
    .RN(net347),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.a[11] ),
    .QN(_20506_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[12]$_DFF_PN0_  (.D(_00355_),
    .RN(net347),
    .CK(clknet_leaf_77_clk),
    .Q(\g_reduce0[10].adder.a[12] ),
    .QN(_20503_));
 DFFR_X1 \g_row[2].g_col[2].mult.x[13]$_DFF_PN0_  (.D(_00356_),
    .RN(net347),
    .CK(clknet_leaf_77_clk),
    .Q(\g_reduce0[10].adder.a[13] ),
    .QN(_20500_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[14]$_DFF_PN0_  (.D(_00357_),
    .RN(net347),
    .CK(clknet_leaf_77_clk),
    .Q(\g_reduce0[10].adder.a[14] ),
    .QN(_20542_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[15]$_DFF_PN0_  (.D(\g_row[2].g_col[2].mult.sign ),
    .RN(net346),
    .CK(clknet_leaf_111_clk),
    .Q(\g_reduce0[10].adder.a[15] ),
    .QN(_13838_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[1]$_DFF_PN0_  (.D(_00358_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.a[1] ),
    .QN(_20536_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[2]$_DFF_PN0_  (.D(_00359_),
    .RN(net346),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.a[2] ),
    .QN(_20533_));
 DFFR_X1 \g_row[2].g_col[2].mult.x[3]$_DFF_PN0_  (.D(_00360_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.a[3] ),
    .QN(_20530_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[4]$_DFF_PN0_  (.D(_00361_),
    .RN(net346),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.a[4] ),
    .QN(_20527_));
 DFFR_X1 \g_row[2].g_col[2].mult.x[5]$_DFF_PN0_  (.D(_00362_),
    .RN(net347),
    .CK(clknet_leaf_71_clk),
    .Q(\g_reduce0[10].adder.a[5] ),
    .QN(_20524_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[6]$_DFF_PN0_  (.D(_00363_),
    .RN(net346),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.a[6] ),
    .QN(_20521_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[7]$_DFF_PN0_  (.D(_00364_),
    .RN(net346),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.a[7] ),
    .QN(_20518_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[8]$_DFF_PN0_  (.D(_00365_),
    .RN(net346),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.a[8] ),
    .QN(_20515_));
 DFFR_X2 \g_row[2].g_col[2].mult.x[9]$_DFF_PN0_  (.D(_00366_),
    .RN(net347),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.a[9] ),
    .QN(_20512_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.expa[0]$_DFF_PN0_  (.D(net85),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_row[2].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14411_));
 DFFR_X2 \g_row[2].g_col[3].mult.stage1.expa[1]$_DFF_PN0_  (.D(net86),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_row[2].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14415_));
 DFFR_X2 \g_row[2].g_col[3].mult.stage1.expa[2]$_DFF_PN0_  (.D(net87),
    .RN(net348),
    .CK(clknet_leaf_124_clk),
    .Q(\g_row[2].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13839_));
 DFFR_X2 \g_row[2].g_col[3].mult.stage1.expa[3]$_DFF_PN0_  (.D(net88),
    .RN(net348),
    .CK(clknet_leaf_124_clk),
    .Q(\g_row[2].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13840_));
 DFFR_X2 \g_row[2].g_col[3].mult.stage1.expa[4]$_DFF_PN0_  (.D(net90),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[2].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13841_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.sign$_DFF_PN0_  (.D(_00383_),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_row[2].g_col[3].mult.sign ),
    .QN(_13842_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[0] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[0] ),
    .QN(_13843_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[10] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[10] ),
    .QN(_13844_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[11] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[11] ),
    .QN(_13845_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[12] ),
    .RN(net349),
    .CK(clknet_leaf_147_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[12] ),
    .QN(_13846_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[13] ),
    .RN(net350),
    .CK(clknet_leaf_165_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[13] ),
    .QN(_13847_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[14] ),
    .RN(net350),
    .CK(clknet_leaf_165_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[14] ),
    .QN(_13848_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[15] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[15] ),
    .QN(_13849_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[16] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[16] ),
    .QN(_13850_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[17] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[17] ),
    .QN(_13851_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[18] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[18] ),
    .QN(_13852_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[19] ),
    .RN(net350),
    .CK(clknet_leaf_160_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[19] ),
    .QN(_13853_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[1] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[1] ),
    .QN(_13854_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[2] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[2] ),
    .QN(_14406_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[3] ),
    .RN(net349),
    .CK(clknet_leaf_149_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[3] ),
    .QN(_13855_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[4] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[4] ),
    .QN(_13856_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[5] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[5] ),
    .QN(_13857_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[6] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[6] ),
    .QN(_13858_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[7] ),
    .RN(net349),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[7] ),
    .QN(_13859_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[8] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[8] ),
    .QN(_13860_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t1[9] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.a[9] ),
    .QN(_13861_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[10] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[10] ),
    .QN(_13862_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[11] ),
    .RN(net349),
    .CK(clknet_leaf_147_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[11] ),
    .QN(_13863_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[12] ),
    .RN(net350),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[12] ),
    .QN(_13864_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[13] ),
    .RN(net350),
    .CK(clknet_leaf_165_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[13] ),
    .QN(_13865_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[14] ),
    .RN(net350),
    .CK(clknet_leaf_165_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[14] ),
    .QN(_13866_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[15] ),
    .RN(net350),
    .CK(clknet_leaf_165_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[15] ),
    .QN(_13867_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[16] ),
    .RN(net350),
    .CK(clknet_leaf_147_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[16] ),
    .QN(_13868_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[17] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[17] ),
    .QN(_13869_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[18] ),
    .RN(net350),
    .CK(clknet_leaf_164_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[18] ),
    .QN(_13870_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[19] ),
    .RN(net350),
    .CK(clknet_leaf_160_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[19] ),
    .QN(_13871_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[1] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[1] ),
    .QN(_13872_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[20] ),
    .RN(net350),
    .CK(clknet_leaf_159_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[20] ),
    .QN(_13873_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[2] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[2] ),
    .QN(_14407_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[3] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[3] ),
    .QN(_13874_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[4] ),
    .RN(net349),
    .CK(clknet_leaf_149_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[4] ),
    .QN(_13875_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[5] ),
    .RN(net349),
    .CK(clknet_leaf_148_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[5] ),
    .QN(_13876_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[6] ),
    .RN(net349),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[6] ),
    .QN(_13877_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[7] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[7] ),
    .QN(_13878_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[8] ),
    .RN(net349),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[8] ),
    .QN(_13879_));
 DFFR_X1 \g_row[2].g_col[3].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.stage1.dadda.t2[9] ),
    .RN(net349),
    .CK(clknet_leaf_146_clk),
    .Q(\g_row[2].g_col[3].mult.adder.b[9] ),
    .QN(_13880_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[0]$_DFF_PN0_  (.D(_00368_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.b[0] ),
    .QN(_00463_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[10]$_DFF_PN0_  (.D(_00369_),
    .RN(net349),
    .CK(clknet_leaf_113_clk),
    .Q(\g_reduce0[10].adder.b[10] ),
    .QN(_20509_));
 DFFR_X2 \g_row[2].g_col[3].mult.x[11]$_DFF_PN0_  (.D(_00370_),
    .RN(net347),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[10].adder.b[11] ),
    .QN(_00467_));
 DFFR_X2 \g_row[2].g_col[3].mult.x[12]$_DFF_PN0_  (.D(_00371_),
    .RN(net347),
    .CK(clknet_leaf_73_clk),
    .Q(\g_reduce0[10].adder.b[12] ),
    .QN(_00472_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[13]$_DFF_PN0_  (.D(_00372_),
    .RN(net347),
    .CK(clknet_leaf_112_clk),
    .Q(\g_reduce0[10].adder.b[13] ),
    .QN(_00475_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[14]$_DFF_PN0_  (.D(_00373_),
    .RN(net349),
    .CK(clknet_leaf_113_clk),
    .Q(\g_reduce0[10].adder.b[14] ),
    .QN(_13881_));
 DFFR_X2 \g_row[2].g_col[3].mult.x[15]$_DFF_PN0_  (.D(\g_row[2].g_col[3].mult.sign ),
    .RN(net349),
    .CK(clknet_leaf_110_clk),
    .Q(\g_reduce0[10].adder.b[15] ),
    .QN(_13882_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[1]$_DFF_PN0_  (.D(_00374_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.b[1] ),
    .QN(_00462_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[2]$_DFF_PN0_  (.D(_00375_),
    .RN(net347),
    .CK(clknet_leaf_72_clk),
    .Q(\g_reduce0[10].adder.b[2] ),
    .QN(_00466_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[3]$_DFF_PN0_  (.D(_00376_),
    .RN(net347),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[10].adder.b[3] ),
    .QN(_00465_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[4]$_DFF_PN0_  (.D(_00377_),
    .RN(net347),
    .CK(clknet_leaf_115_clk),
    .Q(\g_reduce0[10].adder.b[4] ),
    .QN(_00469_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[5]$_DFF_PN0_  (.D(_00378_),
    .RN(net347),
    .CK(clknet_leaf_115_clk),
    .Q(\g_reduce0[10].adder.b[5] ),
    .QN(_00468_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[6]$_DFF_PN0_  (.D(_00379_),
    .RN(net347),
    .CK(clknet_leaf_115_clk),
    .Q(\g_reduce0[10].adder.b[6] ),
    .QN(_00471_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[7]$_DFF_PN0_  (.D(_00380_),
    .RN(net347),
    .CK(clknet_leaf_115_clk),
    .Q(\g_reduce0[10].adder.b[7] ),
    .QN(_00470_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[8]$_DFF_PN0_  (.D(_00381_),
    .RN(net347),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[10].adder.b[8] ),
    .QN(_00474_));
 DFFR_X1 \g_row[2].g_col[3].mult.x[9]$_DFF_PN0_  (.D(_00382_),
    .RN(net349),
    .CK(clknet_leaf_114_clk),
    .Q(\g_reduce0[10].adder.b[9] ),
    .QN(_00473_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.expa[0]$_DFF_PN0_  (.D(net102),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_row[3].g_col[0].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14428_));
 DFFR_X2 \g_row[3].g_col[0].mult.stage1.expa[1]$_DFF_PN0_  (.D(net103),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_row[3].g_col[0].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14432_));
 DFFR_X2 \g_row[3].g_col[0].mult.stage1.expa[2]$_DFF_PN0_  (.D(net104),
    .RN(net350),
    .CK(clknet_leaf_170_clk),
    .Q(\g_row[3].g_col[0].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13883_));
 DFFR_X2 \g_row[3].g_col[0].mult.stage1.expa[3]$_DFF_PN0_  (.D(net105),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[3].g_col[0].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13884_));
 DFFR_X2 \g_row[3].g_col[0].mult.stage1.expa[4]$_DFF_PN0_  (.D(net106),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[3].g_col[0].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13885_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.sign$_DFF_PN0_  (.D(_00399_),
    .RN(net350),
    .CK(clknet_leaf_168_clk),
    .Q(\g_row[3].g_col[0].mult.sign ),
    .QN(_13886_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[0] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[0] ),
    .QN(_13887_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[10] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[10] ),
    .QN(_13888_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[11] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[11] ),
    .QN(_13889_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[12] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[12] ),
    .QN(_13890_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[13] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[13] ),
    .QN(_13891_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[14] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[14] ),
    .QN(_13892_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[15] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[15] ),
    .QN(_13893_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[16] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[16] ),
    .QN(_13894_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[17] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[17] ),
    .QN(_13895_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[18] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[18] ),
    .QN(_13896_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[19] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[19] ),
    .QN(_13897_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[1] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[1] ),
    .QN(_13898_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[2] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[2] ),
    .QN(_14423_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[3] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[3] ),
    .QN(_13899_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[4] ),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[4] ),
    .QN(_13900_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[5] ),
    .RN(net351),
    .CK(clknet_leaf_37_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[5] ),
    .QN(_13901_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[6] ),
    .RN(net351),
    .CK(clknet_leaf_37_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[6] ),
    .QN(_13902_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[7] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[7] ),
    .QN(_13903_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[8] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[8] ),
    .QN(_13904_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t1[9] ),
    .RN(net351),
    .CK(clknet_leaf_36_clk),
    .Q(\g_row[3].g_col[0].mult.adder.a[9] ),
    .QN(_13905_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[10] ),
    .RN(net351),
    .CK(clknet_leaf_36_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[10] ),
    .QN(_13906_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[11] ),
    .RN(net351),
    .CK(clknet_leaf_38_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[11] ),
    .QN(_13907_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[12] ),
    .RN(net351),
    .CK(clknet_leaf_36_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[12] ),
    .QN(_13908_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[13] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[13] ),
    .QN(_13909_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[14] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[14] ),
    .QN(_13910_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[15] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[15] ),
    .QN(_13911_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[16] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[16] ),
    .QN(_13912_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[17] ),
    .RN(net351),
    .CK(clknet_leaf_11_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[17] ),
    .QN(_13913_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[18] ),
    .RN(net351),
    .CK(clknet_leaf_8_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[18] ),
    .QN(_13914_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[19] ),
    .RN(net351),
    .CK(clknet_leaf_9_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[19] ),
    .QN(_13915_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[1] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[1] ),
    .QN(_13916_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[20] ),
    .RN(net347),
    .CK(clknet_leaf_12_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[20] ),
    .QN(_13917_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[2] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[2] ),
    .QN(_14424_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[3] ),
    .RN(net351),
    .CK(clknet_leaf_31_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[3] ),
    .QN(_13918_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[4] ),
    .RN(net351),
    .CK(clknet_leaf_32_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[4] ),
    .QN(_13919_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[5] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[5] ),
    .QN(_13920_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[6] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[6] ),
    .QN(_13921_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[7] ),
    .RN(net351),
    .CK(clknet_leaf_35_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[7] ),
    .QN(_13922_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[8] ),
    .RN(net351),
    .CK(clknet_leaf_36_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[8] ),
    .QN(_13923_));
 DFFR_X1 \g_row[3].g_col[0].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.stage1.dadda.t2[9] ),
    .RN(net351),
    .CK(clknet_leaf_36_clk),
    .Q(\g_row[3].g_col[0].mult.adder.b[9] ),
    .QN(_13924_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[0]$_DFF_PN0_  (.D(_00384_),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_reduce0[12].adder.a[0] ),
    .QN(_00478_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[10]$_DFF_PN0_  (.D(_00385_),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_reduce0[12].adder.a[10] ),
    .QN(_13925_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[11]$_DFF_PN0_  (.D(_00386_),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_reduce0[12].adder.a[11] ),
    .QN(_21124_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[12]$_DFF_PN0_  (.D(_00387_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.a[12] ),
    .QN(_21121_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[13]$_DFF_PN0_  (.D(_00388_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.a[13] ),
    .QN(_21118_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[14]$_DFF_PN0_  (.D(_00389_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.a[14] ),
    .QN(_21160_));
 DFFR_X2 \g_row[3].g_col[0].mult.x[15]$_DFF_PN0_  (.D(\g_row[3].g_col[0].mult.sign ),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_reduce0[12].adder.a[15] ),
    .QN(_13926_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[1]$_DFF_PN0_  (.D(_00390_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.a[1] ),
    .QN(_21154_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[2]$_DFF_PN0_  (.D(_00391_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.a[2] ),
    .QN(_21151_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[3]$_DFF_PN0_  (.D(_00392_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.a[3] ),
    .QN(_21148_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[4]$_DFF_PN0_  (.D(_00393_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.a[4] ),
    .QN(_21145_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[5]$_DFF_PN0_  (.D(_00394_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.a[5] ),
    .QN(_21142_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[6]$_DFF_PN0_  (.D(_00395_),
    .RN(net276),
    .CK(clknet_leaf_20_clk),
    .Q(\g_reduce0[12].adder.a[6] ),
    .QN(_21139_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[7]$_DFF_PN0_  (.D(_00396_),
    .RN(net276),
    .CK(clknet_leaf_20_clk),
    .Q(\g_reduce0[12].adder.a[7] ),
    .QN(_21136_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[8]$_DFF_PN0_  (.D(_00397_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.a[8] ),
    .QN(_21133_));
 DFFR_X1 \g_row[3].g_col[0].mult.x[9]$_DFF_PN0_  (.D(_00398_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.a[9] ),
    .QN(_21130_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.expa[0]$_DFF_PN0_  (.D(net118),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_row[3].g_col[1].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14445_));
 DFFR_X2 \g_row[3].g_col[1].mult.stage1.expa[1]$_DFF_PN0_  (.D(net119),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_row[3].g_col[1].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14449_));
 DFFR_X2 \g_row[3].g_col[1].mult.stage1.expa[2]$_DFF_PN0_  (.D(net121),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[3].g_col[1].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13927_));
 DFFR_X2 \g_row[3].g_col[1].mult.stage1.expa[3]$_DFF_PN0_  (.D(net122),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[3].g_col[1].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13928_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.expa[4]$_DFF_PN0_  (.D(net123),
    .RN(net350),
    .CK(clknet_leaf_169_clk),
    .Q(\g_row[3].g_col[1].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13929_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.sign$_DFF_PN0_  (.D(_00415_),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_row[3].g_col[1].mult.sign ),
    .QN(_13930_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[0] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[0] ),
    .QN(_13931_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[10] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[10] ),
    .QN(_13932_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[11] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[11] ),
    .QN(_13933_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[12] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[12] ),
    .QN(_13934_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[13] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[13] ),
    .QN(_13935_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[14] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[14] ),
    .QN(_13936_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[15] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[15] ),
    .QN(_13937_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[16] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[16] ),
    .QN(_13938_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[17] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[17] ),
    .QN(_13939_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[18] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[18] ),
    .QN(_13940_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[19] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[19] ),
    .QN(_13941_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[1] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[1] ),
    .QN(_13942_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[2] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[2] ),
    .QN(_14440_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[3] ),
    .RN(net276),
    .CK(clknet_leaf_174_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[3] ),
    .QN(_13943_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[4] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[4] ),
    .QN(_13944_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[5] ),
    .RN(net276),
    .CK(clknet_leaf_176_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[5] ),
    .QN(_13945_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[6] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[6] ),
    .QN(_13946_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[7] ),
    .RN(net276),
    .CK(clknet_leaf_3_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[7] ),
    .QN(_13947_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[8] ),
    .RN(net276),
    .CK(clknet_leaf_3_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[8] ),
    .QN(_13948_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t1[9] ),
    .RN(net351),
    .CK(clknet_leaf_3_clk),
    .Q(\g_row[3].g_col[1].mult.adder.a[9] ),
    .QN(_13949_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[10] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[10] ),
    .QN(_13950_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[11] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[11] ),
    .QN(_13951_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[12] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[12] ),
    .QN(_13952_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[13] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[13] ),
    .QN(_13953_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[14] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[14] ),
    .QN(_13954_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[15] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[15] ),
    .QN(_13955_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[16] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[16] ),
    .QN(_13956_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[17] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[17] ),
    .QN(_13957_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[18] ),
    .RN(net351),
    .CK(clknet_leaf_0_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[18] ),
    .QN(_13958_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[19] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[19] ),
    .QN(_13959_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[1] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[1] ),
    .QN(_13960_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[20] ),
    .RN(net351),
    .CK(clknet_leaf_1_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[20] ),
    .QN(_13961_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[2] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[2] ),
    .QN(_14441_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[3] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[3] ),
    .QN(_13962_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[4] ),
    .RN(net276),
    .CK(clknet_leaf_175_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[4] ),
    .QN(_13963_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[5] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[5] ),
    .QN(_13964_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[6] ),
    .RN(net276),
    .CK(clknet_leaf_177_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[6] ),
    .QN(_13965_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[7] ),
    .RN(net276),
    .CK(clknet_leaf_3_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[7] ),
    .QN(_13966_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[8] ),
    .RN(net276),
    .CK(clknet_leaf_3_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[8] ),
    .QN(_13967_));
 DFFR_X1 \g_row[3].g_col[1].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.stage1.dadda.t2[9] ),
    .RN(net351),
    .CK(clknet_leaf_2_clk),
    .Q(\g_row[3].g_col[1].mult.adder.b[9] ),
    .QN(_13968_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[0]$_DFF_PN0_  (.D(_00400_),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_reduce0[12].adder.b[0] ),
    .QN(_00477_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[10]$_DFF_PN0_  (.D(_00401_),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_reduce0[12].adder.b[10] ),
    .QN(_21127_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[11]$_DFF_PN0_  (.D(_00402_),
    .RN(net276),
    .CK(clknet_leaf_162_clk),
    .Q(\g_reduce0[12].adder.b[11] ),
    .QN(_00481_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[12]$_DFF_PN0_  (.D(_00403_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.b[12] ),
    .QN(_00486_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[13]$_DFF_PN0_  (.D(_00404_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.b[13] ),
    .QN(_00489_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[14]$_DFF_PN0_  (.D(_00405_),
    .RN(net276),
    .CK(clknet_leaf_163_clk),
    .Q(\g_reduce0[12].adder.b[14] ),
    .QN(_13969_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[15]$_DFF_PN0_  (.D(\g_row[3].g_col[1].mult.sign ),
    .RN(net350),
    .CK(clknet_leaf_167_clk),
    .Q(\g_reduce0[12].adder.b[15] ),
    .QN(_13970_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[1]$_DFF_PN0_  (.D(_00406_),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_reduce0[12].adder.b[1] ),
    .QN(_00476_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[2]$_DFF_PN0_  (.D(_00407_),
    .RN(net276),
    .CK(clknet_leaf_161_clk),
    .Q(\g_reduce0[12].adder.b[2] ),
    .QN(_00480_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[3]$_DFF_PN0_  (.D(_00408_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.b[3] ),
    .QN(_00479_));
 DFFR_X1 \g_row[3].g_col[1].mult.x[4]$_DFF_PN0_  (.D(_00409_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.b[4] ),
    .QN(_00483_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[5]$_DFF_PN0_  (.D(_00410_),
    .RN(net276),
    .CK(clknet_leaf_18_clk),
    .Q(\g_reduce0[12].adder.b[5] ),
    .QN(_00482_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[6]$_DFF_PN0_  (.D(_00411_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.b[6] ),
    .QN(_00485_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[7]$_DFF_PN0_  (.D(_00412_),
    .RN(net276),
    .CK(clknet_leaf_20_clk),
    .Q(\g_reduce0[12].adder.b[7] ),
    .QN(_00484_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[8]$_DFF_PN0_  (.D(_00413_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.b[8] ),
    .QN(_00488_));
 DFFR_X2 \g_row[3].g_col[1].mult.x[9]$_DFF_PN0_  (.D(_00414_),
    .RN(net276),
    .CK(clknet_leaf_19_clk),
    .Q(\g_reduce0[12].adder.b[9] ),
    .QN(_00487_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.expa[0]$_DFF_PN0_  (.D(net135),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[3].g_col[2].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14462_));
 DFFR_X2 \g_row[3].g_col[2].mult.stage1.expa[1]$_DFF_PN0_  (.D(net136),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[3].g_col[2].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14467_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.expa[2]$_DFF_PN0_  (.D(net137),
    .RN(net346),
    .CK(clknet_leaf_78_clk),
    .Q(\g_row[3].g_col[2].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_13971_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.expa[3]$_DFF_PN0_  (.D(net138),
    .RN(net346),
    .CK(clknet_leaf_93_clk),
    .Q(\g_row[3].g_col[2].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_13972_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.expa[4]$_DFF_PN0_  (.D(net139),
    .RN(net346),
    .CK(clknet_leaf_93_clk),
    .Q(\g_row[3].g_col[2].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_13973_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.sign$_DFF_PN0_  (.D(_00431_),
    .RN(net346),
    .CK(clknet_leaf_97_clk),
    .Q(\g_row[3].g_col[2].mult.sign ),
    .QN(_13974_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[0] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[0] ),
    .QN(_13975_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[10] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[10] ),
    .QN(_13976_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[11] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[11] ),
    .QN(_13977_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[12] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[12] ),
    .QN(_13978_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[13] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[13] ),
    .QN(_13979_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[14] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[14] ),
    .QN(_13980_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[15] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[15] ),
    .QN(_13981_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[16] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[16] ),
    .QN(_13982_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[17] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[17] ),
    .QN(_13983_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[18] ),
    .RN(net345),
    .CK(clknet_leaf_68_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[18] ),
    .QN(_13984_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[19] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[19] ),
    .QN(_13985_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[1] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[1] ),
    .QN(_13986_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[2] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[2] ),
    .QN(_14457_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[3] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[3] ),
    .QN(_13987_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[4] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[4] ),
    .QN(_13988_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[5] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[5] ),
    .QN(_13989_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[6] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[6] ),
    .QN(_13990_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[7] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[7] ),
    .QN(_13991_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[8] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[8] ),
    .QN(_13992_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t1[9] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.a[9] ),
    .QN(_13993_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[10] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[10] ),
    .QN(_13994_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[11] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[11] ),
    .QN(_13995_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[12] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[12] ),
    .QN(_13996_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[13] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[13] ),
    .QN(_13997_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[14] ),
    .RN(net345),
    .CK(clknet_leaf_57_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[14] ),
    .QN(_13998_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[15] ),
    .RN(net345),
    .CK(clknet_leaf_56_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[15] ),
    .QN(_13999_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[16] ),
    .RN(net345),
    .CK(clknet_leaf_67_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[16] ),
    .QN(_14000_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[17] ),
    .RN(net345),
    .CK(clknet_leaf_68_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[17] ),
    .QN(_14001_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[18] ),
    .RN(net345),
    .CK(clknet_leaf_68_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[18] ),
    .QN(_14002_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[19] ),
    .RN(net345),
    .CK(clknet_leaf_68_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[19] ),
    .QN(_14003_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[1] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[1] ),
    .QN(_14004_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[20] ),
    .RN(net345),
    .CK(clknet_leaf_68_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[20] ),
    .QN(_14005_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[2] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[2] ),
    .QN(_14458_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[3] ),
    .RN(net345),
    .CK(clknet_leaf_64_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[3] ),
    .QN(_14006_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[4] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[4] ),
    .QN(_14007_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[5] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[5] ),
    .QN(_14008_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[6] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[6] ),
    .QN(_14009_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[7] ),
    .RN(net345),
    .CK(clknet_leaf_65_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[7] ),
    .QN(_14010_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[8] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[8] ),
    .QN(_14011_));
 DFFR_X1 \g_row[3].g_col[2].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.stage1.dadda.t2[9] ),
    .RN(net345),
    .CK(clknet_leaf_66_clk),
    .Q(\g_row[3].g_col[2].mult.adder.b[9] ),
    .QN(_14012_));
 DFFR_X2 \g_row[3].g_col[2].mult.x[0]$_DFF_PN0_  (.D(_00416_),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_reduce0[14].adder.a[0] ),
    .QN(_21298_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[10]$_DFF_PN0_  (.D(_00417_),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_reduce0[14].adder.a[10] ),
    .QN(_21301_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[11]$_DFF_PN0_  (.D(_00418_),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_reduce0[14].adder.a[11] ),
    .QN(_00495_));
 DFFR_X2 \g_row[3].g_col[2].mult.x[12]$_DFF_PN0_  (.D(_00419_),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_reduce0[14].adder.a[12] ),
    .QN(_00500_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[13]$_DFF_PN0_  (.D(_00420_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.a[13] ),
    .QN(_00503_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[14]$_DFF_PN0_  (.D(_00421_),
    .RN(net349),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[14].adder.a[14] ),
    .QN(_14013_));
 DFFR_X2 \g_row[3].g_col[2].mult.x[15]$_DFF_PN0_  (.D(\g_row[3].g_col[2].mult.sign ),
    .RN(net349),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[14].adder.a[15] ),
    .QN(_14014_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[1]$_DFF_PN0_  (.D(_00422_),
    .RN(net348),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[14].adder.a[1] ),
    .QN(_00490_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[2]$_DFF_PN0_  (.D(_00423_),
    .RN(net348),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[14].adder.a[2] ),
    .QN(_00494_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[3]$_DFF_PN0_  (.D(_00424_),
    .RN(net348),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[14].adder.a[3] ),
    .QN(_00493_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[4]$_DFF_PN0_  (.D(_00425_),
    .RN(net348),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[14].adder.a[4] ),
    .QN(_00497_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[5]$_DFF_PN0_  (.D(_00426_),
    .RN(net348),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[14].adder.a[5] ),
    .QN(_00496_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[6]$_DFF_PN0_  (.D(_00427_),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_reduce0[14].adder.a[6] ),
    .QN(_00499_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[7]$_DFF_PN0_  (.D(_00428_),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_reduce0[14].adder.a[7] ),
    .QN(_00498_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[8]$_DFF_PN0_  (.D(_00429_),
    .RN(net348),
    .CK(clknet_leaf_108_clk),
    .Q(\g_reduce0[14].adder.a[8] ),
    .QN(_00502_));
 DFFR_X1 \g_row[3].g_col[2].mult.x[9]$_DFF_PN0_  (.D(_00430_),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_reduce0[14].adder.a[9] ),
    .QN(_00501_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.expa[0]$_DFF_PN0_  (.D(net150),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_row[3].g_col[3].mult.expAdder.g_intermediate[0].fa.a ),
    .QN(_14480_));
 DFFR_X2 \g_row[3].g_col[3].mult.stage1.expa[1]$_DFF_PN0_  (.D(net151),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_row[3].g_col[3].mult.expAdder.g_intermediate[1].fa.a ),
    .QN(_14484_));
 DFFR_X2 \g_row[3].g_col[3].mult.stage1.expa[2]$_DFF_PN0_  (.D(net152),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[3].g_col[3].mult.expAdder.g_intermediate[2].fa.a ),
    .QN(_14015_));
 DFFR_X2 \g_row[3].g_col[3].mult.stage1.expa[3]$_DFF_PN0_  (.D(net153),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[3].g_col[3].mult.expAdder.g_intermediate[3].fa.a ),
    .QN(_14016_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.expa[4]$_DFF_PN0_  (.D(net154),
    .RN(net348),
    .CK(clknet_leaf_123_clk),
    .Q(\g_row[3].g_col[3].mult.expAdder.g_intermediate[4].fa.a ),
    .QN(_14017_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.sign$_DFF_PN0_  (.D(_00447_),
    .RN(net349),
    .CK(clknet_leaf_108_clk),
    .Q(\g_row[3].g_col[3].mult.sign ),
    .QN(_14018_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[0]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[0] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[0] ),
    .QN(_14019_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[10]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[10] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[10] ),
    .QN(_14020_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[11]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[11] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[11] ),
    .QN(_14021_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[12]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[12] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[12] ),
    .QN(_14022_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[13]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[13] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[13] ),
    .QN(_14023_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[14]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[14] ),
    .RN(net349),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[14] ),
    .QN(_14024_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[15]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[15] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[15] ),
    .QN(_14025_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[16]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[16] ),
    .RN(net348),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[16] ),
    .QN(_14026_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[17]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[17] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[17] ),
    .QN(_14027_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[18]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[18] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[18] ),
    .QN(_14028_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[19]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[19] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[19] ),
    .QN(_14029_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[1]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[1] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[1] ),
    .QN(_14030_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[2]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[2] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[2] ),
    .QN(_14475_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[3]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[3] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[3] ),
    .QN(_14031_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[4]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[4] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[4] ),
    .QN(_14032_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[5]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[5] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[5] ),
    .QN(_14033_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[6]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[6] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[6] ),
    .QN(_14034_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[7]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[7] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[7] ),
    .QN(_14035_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[8]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[8] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[8] ),
    .QN(_14036_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t1[9]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t1[9] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.a[9] ),
    .QN(_14037_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[10]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[10] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[10] ),
    .QN(_14038_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[11]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[11] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[11] ),
    .QN(_14039_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[12]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[12] ),
    .RN(net349),
    .CK(clknet_leaf_142_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[12] ),
    .QN(_14040_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[13]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[13] ),
    .RN(net349),
    .CK(clknet_leaf_145_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[13] ),
    .QN(_14041_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[14]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[14] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[14] ),
    .QN(_14042_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[15]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[15] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[15] ),
    .QN(_14043_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[16]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[16] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[16] ),
    .QN(_14044_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[17]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[17] ),
    .RN(net349),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[17] ),
    .QN(_14045_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[18]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[18] ),
    .RN(net348),
    .CK(clknet_leaf_141_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[18] ),
    .QN(_14046_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[19]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[19] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[19] ),
    .QN(_14047_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[1]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[1] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[1] ),
    .QN(_14048_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[20]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[20] ),
    .RN(net348),
    .CK(clknet_leaf_140_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[20] ),
    .QN(_14049_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[2]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[2] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[2] ),
    .QN(_14476_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[3]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[3] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[3] ),
    .QN(_14050_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[4]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[4] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[4] ),
    .QN(_14051_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[5]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[5] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[5] ),
    .QN(_14052_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[6]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[6] ),
    .RN(net349),
    .CK(clknet_leaf_134_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[6] ),
    .QN(_14053_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[7]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[7] ),
    .RN(net349),
    .CK(clknet_leaf_144_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[7] ),
    .QN(_14054_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[8]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[8] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[8] ),
    .QN(_14055_));
 DFFR_X1 \g_row[3].g_col[3].mult.stage1.t2[9]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.stage1.dadda.t2[9] ),
    .RN(net349),
    .CK(clknet_leaf_143_clk),
    .Q(\g_row[3].g_col[3].mult.adder.b[9] ),
    .QN(_14056_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[0]$_DFF_PN0_  (.D(_00432_),
    .RN(net348),
    .CK(clknet_leaf_107_clk),
    .Q(\g_reduce0[14].adder.b[0] ),
    .QN(_00491_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[10]$_DFF_PN0_  (.D(_00433_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.b[10] ),
    .QN(_00492_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[11]$_DFF_PN0_  (.D(_00434_),
    .RN(net348),
    .CK(clknet_leaf_106_clk),
    .Q(\g_reduce0[14].adder.b[11] ),
    .QN(_21268_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[12]$_DFF_PN0_  (.D(_00435_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[14].adder.b[12] ),
    .QN(_21265_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[13]$_DFF_PN0_  (.D(_00436_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[14].adder.b[13] ),
    .QN(_21262_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[14]$_DFF_PN0_  (.D(_00437_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[14].adder.b[14] ),
    .QN(_21307_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[15]$_DFF_PN0_  (.D(\g_row[3].g_col[3].mult.sign ),
    .RN(net349),
    .CK(clknet_leaf_109_clk),
    .Q(\g_reduce0[14].adder.b[15] ),
    .QN(_14057_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[1]$_DFF_PN0_  (.D(_00438_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.b[1] ),
    .QN(_21295_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[2]$_DFF_PN0_  (.D(_00439_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.b[2] ),
    .QN(_21292_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[3]$_DFF_PN0_  (.D(_00440_),
    .RN(net348),
    .CK(clknet_leaf_122_clk),
    .Q(\g_reduce0[14].adder.b[3] ),
    .QN(_21289_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[4]$_DFF_PN0_  (.D(_00441_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.b[4] ),
    .QN(_21286_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[5]$_DFF_PN0_  (.D(_00442_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.b[5] ),
    .QN(_21283_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[6]$_DFF_PN0_  (.D(_00443_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.b[6] ),
    .QN(_21280_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[7]$_DFF_PN0_  (.D(_00444_),
    .RN(net348),
    .CK(clknet_leaf_121_clk),
    .Q(\g_reduce0[14].adder.b[7] ),
    .QN(_21277_));
 DFFR_X1 \g_row[3].g_col[3].mult.x[8]$_DFF_PN0_  (.D(_00445_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.b[8] ),
    .QN(_21274_));
 DFFR_X2 \g_row[3].g_col[3].mult.x[9]$_DFF_PN0_  (.D(_00446_),
    .RN(net348),
    .CK(clknet_leaf_120_clk),
    .Q(\g_reduce0[14].adder.b[9] ),
    .QN(_21271_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_387 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 BUF_X1 input2 (.A(a[100]),
    .Z(net2));
 BUF_X1 input3 (.A(a[101]),
    .Z(net3));
 BUF_X1 input4 (.A(a[102]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(a[104]),
    .Z(net5));
 BUF_X1 input6 (.A(a[106]),
    .Z(net6));
 BUF_X1 input7 (.A(a[107]),
    .Z(net7));
 BUF_X1 input8 (.A(a[108]),
    .Z(net8));
 BUF_X1 input9 (.A(a[109]),
    .Z(net9));
 BUF_X1 input10 (.A(a[10]),
    .Z(net10));
 BUF_X1 input11 (.A(a[110]),
    .Z(net11));
 BUF_X1 input12 (.A(a[111]),
    .Z(net12));
 BUF_X1 input13 (.A(a[112]),
    .Z(net13));
 BUF_X1 input14 (.A(a[113]),
    .Z(net14));
 BUF_X1 input15 (.A(a[114]),
    .Z(net15));
 BUF_X1 input16 (.A(a[115]),
    .Z(net16));
 BUF_X1 input17 (.A(a[116]),
    .Z(net17));
 BUF_X1 input18 (.A(a[117]),
    .Z(net18));
 BUF_X2 input19 (.A(a[118]),
    .Z(net19));
 BUF_X1 input20 (.A(a[11]),
    .Z(net20));
 BUF_X2 input21 (.A(a[120]),
    .Z(net21));
 BUF_X1 input22 (.A(a[122]),
    .Z(net22));
 BUF_X1 input23 (.A(a[123]),
    .Z(net23));
 BUF_X1 input24 (.A(a[124]),
    .Z(net24));
 BUF_X1 input25 (.A(a[125]),
    .Z(net25));
 BUF_X1 input26 (.A(a[126]),
    .Z(net26));
 BUF_X1 input27 (.A(a[127]),
    .Z(net27));
 BUF_X1 input28 (.A(a[128]),
    .Z(net28));
 BUF_X1 input29 (.A(a[129]),
    .Z(net29));
 BUF_X1 input30 (.A(a[12]),
    .Z(net30));
 BUF_X1 input31 (.A(a[130]),
    .Z(net31));
 BUF_X1 input32 (.A(a[131]),
    .Z(net32));
 BUF_X1 input33 (.A(a[132]),
    .Z(net33));
 BUF_X1 input34 (.A(a[133]),
    .Z(net34));
 BUF_X1 input35 (.A(a[134]),
    .Z(net35));
 CLKBUF_X2 input36 (.A(a[136]),
    .Z(net36));
 BUF_X1 input37 (.A(a[138]),
    .Z(net37));
 BUF_X1 input38 (.A(a[139]),
    .Z(net38));
 BUF_X1 input39 (.A(a[13]),
    .Z(net39));
 BUF_X1 input40 (.A(a[140]),
    .Z(net40));
 BUF_X1 input41 (.A(a[141]),
    .Z(net41));
 BUF_X1 input42 (.A(a[142]),
    .Z(net42));
 BUF_X1 input43 (.A(a[143]),
    .Z(net43));
 BUF_X1 input44 (.A(a[144]),
    .Z(net44));
 BUF_X1 input45 (.A(a[145]),
    .Z(net45));
 BUF_X1 input46 (.A(a[146]),
    .Z(net46));
 BUF_X1 input47 (.A(a[147]),
    .Z(net47));
 BUF_X1 input48 (.A(a[148]),
    .Z(net48));
 BUF_X1 input49 (.A(a[149]),
    .Z(net49));
 BUF_X1 input50 (.A(a[14]),
    .Z(net50));
 BUF_X1 input51 (.A(a[150]),
    .Z(net51));
 BUF_X1 input52 (.A(a[151]),
    .Z(net52));
 CLKBUF_X2 input53 (.A(a[152]),
    .Z(net53));
 BUF_X1 input54 (.A(a[154]),
    .Z(net54));
 BUF_X1 input55 (.A(a[155]),
    .Z(net55));
 BUF_X1 input56 (.A(a[156]),
    .Z(net56));
 BUF_X1 input57 (.A(a[157]),
    .Z(net57));
 BUF_X1 input58 (.A(a[158]),
    .Z(net58));
 BUF_X1 input59 (.A(a[159]),
    .Z(net59));
 BUF_X1 input60 (.A(a[15]),
    .Z(net60));
 BUF_X1 input61 (.A(a[160]),
    .Z(net61));
 BUF_X1 input62 (.A(a[161]),
    .Z(net62));
 BUF_X1 input63 (.A(a[162]),
    .Z(net63));
 BUF_X1 input64 (.A(a[163]),
    .Z(net64));
 BUF_X1 input65 (.A(a[164]),
    .Z(net65));
 BUF_X1 input66 (.A(a[165]),
    .Z(net66));
 BUF_X1 input67 (.A(a[166]),
    .Z(net67));
 CLKBUF_X2 input68 (.A(a[168]),
    .Z(net68));
 BUF_X1 input69 (.A(a[16]),
    .Z(net69));
 BUF_X1 input70 (.A(a[170]),
    .Z(net70));
 BUF_X1 input71 (.A(a[171]),
    .Z(net71));
 BUF_X1 input72 (.A(a[172]),
    .Z(net72));
 BUF_X1 input73 (.A(a[173]),
    .Z(net73));
 BUF_X1 input74 (.A(a[174]),
    .Z(net74));
 BUF_X1 input75 (.A(a[175]),
    .Z(net75));
 BUF_X1 input76 (.A(a[176]),
    .Z(net76));
 BUF_X1 input77 (.A(a[177]),
    .Z(net77));
 BUF_X1 input78 (.A(a[178]),
    .Z(net78));
 BUF_X1 input79 (.A(a[179]),
    .Z(net79));
 BUF_X1 input80 (.A(a[17]),
    .Z(net80));
 BUF_X1 input81 (.A(a[180]),
    .Z(net81));
 BUF_X1 input82 (.A(a[181]),
    .Z(net82));
 BUF_X1 input83 (.A(a[182]),
    .Z(net83));
 BUF_X2 input84 (.A(a[184]),
    .Z(net84));
 BUF_X1 input85 (.A(a[186]),
    .Z(net85));
 BUF_X1 input86 (.A(a[187]),
    .Z(net86));
 BUF_X1 input87 (.A(a[188]),
    .Z(net87));
 BUF_X1 input88 (.A(a[189]),
    .Z(net88));
 BUF_X1 input89 (.A(a[18]),
    .Z(net89));
 BUF_X1 input90 (.A(a[190]),
    .Z(net90));
 BUF_X1 input91 (.A(a[191]),
    .Z(net91));
 BUF_X1 input92 (.A(a[192]),
    .Z(net92));
 BUF_X1 input93 (.A(a[193]),
    .Z(net93));
 BUF_X1 input94 (.A(a[194]),
    .Z(net94));
 BUF_X1 input95 (.A(a[195]),
    .Z(net95));
 BUF_X1 input96 (.A(a[196]),
    .Z(net96));
 BUF_X1 input97 (.A(a[197]),
    .Z(net97));
 BUF_X1 input98 (.A(a[198]),
    .Z(net98));
 BUF_X1 input99 (.A(a[19]),
    .Z(net99));
 BUF_X1 input100 (.A(a[1]),
    .Z(net100));
 CLKBUF_X2 input101 (.A(a[200]),
    .Z(net101));
 BUF_X1 input102 (.A(a[202]),
    .Z(net102));
 BUF_X1 input103 (.A(a[203]),
    .Z(net103));
 BUF_X1 input104 (.A(a[204]),
    .Z(net104));
 BUF_X1 input105 (.A(a[205]),
    .Z(net105));
 BUF_X1 input106 (.A(a[206]),
    .Z(net106));
 BUF_X1 input107 (.A(a[207]),
    .Z(net107));
 BUF_X1 input108 (.A(a[208]),
    .Z(net108));
 BUF_X1 input109 (.A(a[209]),
    .Z(net109));
 BUF_X1 input110 (.A(a[20]),
    .Z(net110));
 BUF_X1 input111 (.A(a[210]),
    .Z(net111));
 BUF_X1 input112 (.A(a[211]),
    .Z(net112));
 BUF_X1 input113 (.A(a[212]),
    .Z(net113));
 BUF_X1 input114 (.A(a[213]),
    .Z(net114));
 BUF_X1 input115 (.A(a[214]),
    .Z(net115));
 BUF_X1 input116 (.A(a[215]),
    .Z(net116));
 CLKBUF_X2 input117 (.A(a[216]),
    .Z(net117));
 BUF_X1 input118 (.A(a[218]),
    .Z(net118));
 BUF_X1 input119 (.A(a[219]),
    .Z(net119));
 BUF_X1 input120 (.A(a[21]),
    .Z(net120));
 BUF_X1 input121 (.A(a[220]),
    .Z(net121));
 BUF_X1 input122 (.A(a[221]),
    .Z(net122));
 BUF_X1 input123 (.A(a[222]),
    .Z(net123));
 BUF_X1 input124 (.A(a[223]),
    .Z(net124));
 BUF_X1 input125 (.A(a[224]),
    .Z(net125));
 BUF_X1 input126 (.A(a[225]),
    .Z(net126));
 BUF_X1 input127 (.A(a[226]),
    .Z(net127));
 CLKBUF_X2 input128 (.A(a[227]),
    .Z(net128));
 BUF_X2 input129 (.A(a[228]),
    .Z(net129));
 BUF_X2 input130 (.A(a[229]),
    .Z(net130));
 BUF_X1 input131 (.A(a[22]),
    .Z(net131));
 BUF_X2 input132 (.A(a[230]),
    .Z(net132));
 BUF_X2 input133 (.A(a[231]),
    .Z(net133));
 BUF_X2 input134 (.A(a[232]),
    .Z(net134));
 BUF_X1 input135 (.A(a[234]),
    .Z(net135));
 BUF_X1 input136 (.A(a[235]),
    .Z(net136));
 BUF_X1 input137 (.A(a[236]),
    .Z(net137));
 BUF_X1 input138 (.A(a[237]),
    .Z(net138));
 BUF_X1 input139 (.A(a[238]),
    .Z(net139));
 BUF_X1 input140 (.A(a[239]),
    .Z(net140));
 BUF_X1 input141 (.A(a[240]),
    .Z(net141));
 BUF_X1 input142 (.A(a[241]),
    .Z(net142));
 BUF_X1 input143 (.A(a[242]),
    .Z(net143));
 BUF_X1 input144 (.A(a[243]),
    .Z(net144));
 BUF_X1 input145 (.A(a[244]),
    .Z(net145));
 BUF_X1 input146 (.A(a[245]),
    .Z(net146));
 BUF_X1 input147 (.A(a[246]),
    .Z(net147));
 BUF_X2 input148 (.A(a[248]),
    .Z(net148));
 BUF_X2 input149 (.A(a[24]),
    .Z(net149));
 BUF_X1 input150 (.A(a[250]),
    .Z(net150));
 BUF_X1 input151 (.A(a[251]),
    .Z(net151));
 BUF_X1 input152 (.A(a[252]),
    .Z(net152));
 BUF_X1 input153 (.A(a[253]),
    .Z(net153));
 BUF_X1 input154 (.A(a[254]),
    .Z(net154));
 BUF_X1 input155 (.A(a[255]),
    .Z(net155));
 BUF_X1 input156 (.A(a[26]),
    .Z(net156));
 BUF_X1 input157 (.A(a[27]),
    .Z(net157));
 BUF_X1 input158 (.A(a[28]),
    .Z(net158));
 BUF_X1 input159 (.A(a[29]),
    .Z(net159));
 BUF_X1 input160 (.A(a[2]),
    .Z(net160));
 BUF_X1 input161 (.A(a[30]),
    .Z(net161));
 BUF_X1 input162 (.A(a[31]),
    .Z(net162));
 BUF_X1 input163 (.A(a[32]),
    .Z(net163));
 BUF_X1 input164 (.A(a[33]),
    .Z(net164));
 BUF_X1 input165 (.A(a[34]),
    .Z(net165));
 BUF_X1 input166 (.A(a[35]),
    .Z(net166));
 BUF_X1 input167 (.A(a[36]),
    .Z(net167));
 BUF_X1 input168 (.A(a[37]),
    .Z(net168));
 BUF_X1 input169 (.A(a[38]),
    .Z(net169));
 BUF_X1 input170 (.A(a[39]),
    .Z(net170));
 BUF_X1 input171 (.A(a[3]),
    .Z(net171));
 CLKBUF_X3 input172 (.A(a[40]),
    .Z(net172));
 BUF_X1 input173 (.A(a[42]),
    .Z(net173));
 BUF_X1 input174 (.A(a[43]),
    .Z(net174));
 BUF_X1 input175 (.A(a[44]),
    .Z(net175));
 BUF_X1 input176 (.A(a[45]),
    .Z(net176));
 BUF_X1 input177 (.A(a[46]),
    .Z(net177));
 BUF_X1 input178 (.A(a[47]),
    .Z(net178));
 BUF_X1 input179 (.A(a[48]),
    .Z(net179));
 BUF_X1 input180 (.A(a[49]),
    .Z(net180));
 BUF_X1 input181 (.A(a[4]),
    .Z(net181));
 BUF_X1 input182 (.A(a[50]),
    .Z(net182));
 BUF_X1 input183 (.A(a[51]),
    .Z(net183));
 BUF_X1 input184 (.A(a[52]),
    .Z(net184));
 BUF_X1 input185 (.A(a[53]),
    .Z(net185));
 CLKBUF_X2 input186 (.A(a[54]),
    .Z(net186));
 CLKBUF_X3 input187 (.A(a[56]),
    .Z(net187));
 BUF_X1 input188 (.A(a[58]),
    .Z(net188));
 BUF_X1 input189 (.A(a[59]),
    .Z(net189));
 BUF_X1 input190 (.A(a[5]),
    .Z(net190));
 BUF_X1 input191 (.A(a[60]),
    .Z(net191));
 BUF_X1 input192 (.A(a[61]),
    .Z(net192));
 BUF_X1 input193 (.A(a[62]),
    .Z(net193));
 BUF_X1 input194 (.A(a[63]),
    .Z(net194));
 BUF_X1 input195 (.A(a[64]),
    .Z(net195));
 BUF_X1 input196 (.A(a[65]),
    .Z(net196));
 BUF_X1 input197 (.A(a[66]),
    .Z(net197));
 BUF_X1 input198 (.A(a[67]),
    .Z(net198));
 BUF_X1 input199 (.A(a[68]),
    .Z(net199));
 BUF_X1 input200 (.A(a[69]),
    .Z(net200));
 BUF_X1 input201 (.A(a[6]),
    .Z(net201));
 BUF_X1 input202 (.A(a[70]),
    .Z(net202));
 BUF_X1 input203 (.A(a[71]),
    .Z(net203));
 CLKBUF_X2 input204 (.A(a[72]),
    .Z(net204));
 BUF_X1 input205 (.A(a[74]),
    .Z(net205));
 BUF_X1 input206 (.A(a[75]),
    .Z(net206));
 BUF_X1 input207 (.A(a[76]),
    .Z(net207));
 BUF_X1 input208 (.A(a[77]),
    .Z(net208));
 BUF_X1 input209 (.A(a[78]),
    .Z(net209));
 BUF_X1 input210 (.A(a[79]),
    .Z(net210));
 BUF_X1 input211 (.A(a[7]),
    .Z(net211));
 BUF_X1 input212 (.A(a[80]),
    .Z(net212));
 BUF_X1 input213 (.A(a[81]),
    .Z(net213));
 BUF_X1 input214 (.A(a[82]),
    .Z(net214));
 BUF_X1 input215 (.A(a[83]),
    .Z(net215));
 BUF_X1 input216 (.A(a[84]),
    .Z(net216));
 BUF_X1 input217 (.A(a[85]),
    .Z(net217));
 BUF_X1 input218 (.A(a[86]),
    .Z(net218));
 BUF_X1 input219 (.A(a[87]),
    .Z(net219));
 BUF_X2 input220 (.A(a[88]),
    .Z(net220));
 CLKBUF_X2 input221 (.A(a[8]),
    .Z(net221));
 BUF_X1 input222 (.A(a[90]),
    .Z(net222));
 BUF_X1 input223 (.A(a[91]),
    .Z(net223));
 BUF_X1 input224 (.A(a[92]),
    .Z(net224));
 BUF_X1 input225 (.A(a[93]),
    .Z(net225));
 BUF_X1 input226 (.A(a[94]),
    .Z(net226));
 BUF_X1 input227 (.A(a[95]),
    .Z(net227));
 BUF_X1 input228 (.A(a[96]),
    .Z(net228));
 BUF_X1 input229 (.A(a[97]),
    .Z(net229));
 BUF_X1 input230 (.A(a[98]),
    .Z(net230));
 BUF_X1 input231 (.A(a[99]),
    .Z(net231));
 BUF_X1 input232 (.A(b[0]),
    .Z(net232));
 BUF_X1 input233 (.A(b[10]),
    .Z(net233));
 BUF_X1 input234 (.A(b[11]),
    .Z(net234));
 BUF_X1 input235 (.A(b[12]),
    .Z(net235));
 BUF_X1 input236 (.A(b[13]),
    .Z(net236));
 BUF_X1 input237 (.A(b[14]),
    .Z(net237));
 BUF_X1 input238 (.A(b[16]),
    .Z(net238));
 BUF_X1 input239 (.A(b[18]),
    .Z(net239));
 BUF_X1 input240 (.A(b[20]),
    .Z(net240));
 BUF_X4 input241 (.A(b[21]),
    .Z(net241));
 BUF_X4 input242 (.A(b[23]),
    .Z(net242));
 BUF_X1 input243 (.A(b[24]),
    .Z(net243));
 BUF_X1 input244 (.A(b[26]),
    .Z(net244));
 BUF_X1 input245 (.A(b[27]),
    .Z(net245));
 BUF_X1 input246 (.A(b[28]),
    .Z(net246));
 BUF_X1 input247 (.A(b[29]),
    .Z(net247));
 BUF_X1 input248 (.A(b[2]),
    .Z(net248));
 BUF_X1 input249 (.A(b[30]),
    .Z(net249));
 BUF_X1 input250 (.A(b[32]),
    .Z(net250));
 BUF_X1 input251 (.A(b[34]),
    .Z(net251));
 BUF_X4 input252 (.A(b[36]),
    .Z(net252));
 BUF_X1 input253 (.A(b[37]),
    .Z(net253));
 BUF_X4 input254 (.A(b[39]),
    .Z(net254));
 BUF_X1 input255 (.A(b[40]),
    .Z(net255));
 BUF_X1 input256 (.A(b[42]),
    .Z(net256));
 BUF_X1 input257 (.A(b[43]),
    .Z(net257));
 BUF_X1 input258 (.A(b[44]),
    .Z(net258));
 BUF_X1 input259 (.A(b[45]),
    .Z(net259));
 BUF_X1 input260 (.A(b[46]),
    .Z(net260));
 BUF_X1 input261 (.A(b[48]),
    .Z(net261));
 CLKBUF_X3 input262 (.A(b[4]),
    .Z(net262));
 BUF_X1 input263 (.A(b[50]),
    .Z(net263));
 BUF_X4 input264 (.A(b[52]),
    .Z(net264));
 BUF_X1 input265 (.A(b[53]),
    .Z(net265));
 BUF_X4 input266 (.A(b[55]),
    .Z(net266));
 BUF_X1 input267 (.A(b[56]),
    .Z(net267));
 BUF_X1 input268 (.A(b[58]),
    .Z(net268));
 BUF_X1 input269 (.A(b[59]),
    .Z(net269));
 BUF_X1 input270 (.A(b[5]),
    .Z(net270));
 BUF_X1 input271 (.A(b[60]),
    .Z(net271));
 BUF_X1 input272 (.A(b[61]),
    .Z(net272));
 BUF_X1 input273 (.A(b[62]),
    .Z(net273));
 CLKBUF_X3 input274 (.A(b[7]),
    .Z(net274));
 BUF_X1 input275 (.A(b[8]),
    .Z(net275));
 BUF_X1 input276 (.A(rst),
    .Z(net276));
 BUF_X1 output277 (.A(net277),
    .Z(x[0]));
 BUF_X1 output278 (.A(net278),
    .Z(x[10]));
 BUF_X1 output279 (.A(net279),
    .Z(x[11]));
 BUF_X1 output280 (.A(net280),
    .Z(x[12]));
 BUF_X1 output281 (.A(net281),
    .Z(x[13]));
 BUF_X1 output282 (.A(net282),
    .Z(x[14]));
 BUF_X1 output283 (.A(net283),
    .Z(x[15]));
 BUF_X1 output284 (.A(net284),
    .Z(x[16]));
 BUF_X1 output285 (.A(net285),
    .Z(x[17]));
 BUF_X1 output286 (.A(net286),
    .Z(x[18]));
 BUF_X1 output287 (.A(net287),
    .Z(x[19]));
 BUF_X1 output288 (.A(net288),
    .Z(x[1]));
 BUF_X1 output289 (.A(net289),
    .Z(x[20]));
 BUF_X1 output290 (.A(net290),
    .Z(x[21]));
 BUF_X1 output291 (.A(net291),
    .Z(x[22]));
 BUF_X1 output292 (.A(net292),
    .Z(x[23]));
 BUF_X1 output293 (.A(net293),
    .Z(x[24]));
 BUF_X1 output294 (.A(net294),
    .Z(x[25]));
 BUF_X1 output295 (.A(net295),
    .Z(x[26]));
 BUF_X1 output296 (.A(net296),
    .Z(x[27]));
 BUF_X1 output297 (.A(net297),
    .Z(x[28]));
 BUF_X1 output298 (.A(net298),
    .Z(x[29]));
 BUF_X1 output299 (.A(net299),
    .Z(x[2]));
 BUF_X1 output300 (.A(net300),
    .Z(x[30]));
 BUF_X1 output301 (.A(net301),
    .Z(x[31]));
 BUF_X1 output302 (.A(net302),
    .Z(x[32]));
 BUF_X1 output303 (.A(net303),
    .Z(x[33]));
 BUF_X1 output304 (.A(net304),
    .Z(x[34]));
 BUF_X1 output305 (.A(net305),
    .Z(x[35]));
 BUF_X1 output306 (.A(net306),
    .Z(x[36]));
 BUF_X1 output307 (.A(net307),
    .Z(x[37]));
 BUF_X1 output308 (.A(net308),
    .Z(x[38]));
 BUF_X1 output309 (.A(net309),
    .Z(x[39]));
 BUF_X1 output310 (.A(net310),
    .Z(x[3]));
 BUF_X1 output311 (.A(net311),
    .Z(x[40]));
 BUF_X1 output312 (.A(net312),
    .Z(x[41]));
 BUF_X1 output313 (.A(net313),
    .Z(x[42]));
 BUF_X1 output314 (.A(net314),
    .Z(x[43]));
 BUF_X1 output315 (.A(net315),
    .Z(x[44]));
 BUF_X1 output316 (.A(net316),
    .Z(x[45]));
 BUF_X1 output317 (.A(net317),
    .Z(x[46]));
 BUF_X1 output318 (.A(net318),
    .Z(x[47]));
 BUF_X1 output319 (.A(net319),
    .Z(x[48]));
 BUF_X1 output320 (.A(net320),
    .Z(x[49]));
 BUF_X1 output321 (.A(net321),
    .Z(x[4]));
 BUF_X1 output322 (.A(net322),
    .Z(x[50]));
 BUF_X1 output323 (.A(net323),
    .Z(x[51]));
 BUF_X1 output324 (.A(net324),
    .Z(x[52]));
 BUF_X1 output325 (.A(net325),
    .Z(x[53]));
 BUF_X1 output326 (.A(net326),
    .Z(x[54]));
 BUF_X1 output327 (.A(net327),
    .Z(x[55]));
 BUF_X1 output328 (.A(net328),
    .Z(x[56]));
 BUF_X1 output329 (.A(net329),
    .Z(x[57]));
 BUF_X1 output330 (.A(net330),
    .Z(x[58]));
 BUF_X1 output331 (.A(net331),
    .Z(x[59]));
 BUF_X1 output332 (.A(net332),
    .Z(x[5]));
 BUF_X1 output333 (.A(net333),
    .Z(x[60]));
 BUF_X1 output334 (.A(net334),
    .Z(x[61]));
 BUF_X1 output335 (.A(net335),
    .Z(x[62]));
 BUF_X1 output336 (.A(net336),
    .Z(x[63]));
 BUF_X1 output337 (.A(net337),
    .Z(x[6]));
 BUF_X1 output338 (.A(net338),
    .Z(x[7]));
 BUF_X1 output339 (.A(net339),
    .Z(x[8]));
 BUF_X1 output340 (.A(net340),
    .Z(x[9]));
 BUF_X2 max_cap341 (.A(_03064_),
    .Z(net341));
 BUF_X2 max_cap342 (.A(_06368_),
    .Z(net342));
 CLKBUF_X2 max_cap343 (.A(_10419_),
    .Z(net343));
 BUF_X4 wire344 (.A(_10227_),
    .Z(net344));
 BUF_X1 max_length345 (.A(net351),
    .Z(net345));
 BUF_X32 max_length346 (.A(net347),
    .Z(net346));
 BUF_X1 max_length347 (.A(net351),
    .Z(net347));
 BUF_X2 max_length348 (.A(net349),
    .Z(net348));
 BUF_X1 max_length349 (.A(net350),
    .Z(net349));
 BUF_X1 max_length350 (.A(net276),
    .Z(net350));
 BUF_X1 max_length351 (.A(net276),
    .Z(net351));
 BUF_X1 wire352 (.A(a[233]),
    .Z(net352));
 BUF_X1 wire353 (.A(a[121]),
    .Z(net353));
 LOGIC1_X1 \g_row[0].g_col[0].mult.stage1.t1[20]$_DFF_PN0__354  (.Z(net354));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_4_2_0_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_4_10_0_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_4_11_0_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_4_9_0_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_4_14_0_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_leaf_98_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_98_clk));
 CLKBUF_X3 clkbuf_leaf_99_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_99_clk));
 CLKBUF_X3 clkbuf_leaf_100_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_100_clk));
 CLKBUF_X3 clkbuf_leaf_101_clk (.A(clknet_4_15_0_clk),
    .Z(clknet_leaf_101_clk));
 CLKBUF_X3 clkbuf_leaf_102_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_102_clk));
 CLKBUF_X3 clkbuf_leaf_103_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_103_clk));
 CLKBUF_X3 clkbuf_leaf_104_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_104_clk));
 CLKBUF_X3 clkbuf_leaf_105_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_105_clk));
 CLKBUF_X3 clkbuf_leaf_106_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_106_clk));
 CLKBUF_X3 clkbuf_leaf_107_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_107_clk));
 CLKBUF_X3 clkbuf_leaf_108_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_108_clk));
 CLKBUF_X3 clkbuf_leaf_109_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_109_clk));
 CLKBUF_X3 clkbuf_leaf_110_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_110_clk));
 CLKBUF_X3 clkbuf_leaf_111_clk (.A(clknet_4_13_0_clk),
    .Z(clknet_leaf_111_clk));
 CLKBUF_X3 clkbuf_leaf_112_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_112_clk));
 CLKBUF_X3 clkbuf_leaf_113_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_113_clk));
 CLKBUF_X3 clkbuf_leaf_114_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_114_clk));
 CLKBUF_X3 clkbuf_leaf_115_clk (.A(clknet_4_12_0_clk),
    .Z(clknet_leaf_115_clk));
 CLKBUF_X3 clkbuf_leaf_116_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_116_clk));
 CLKBUF_X3 clkbuf_leaf_117_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_117_clk));
 CLKBUF_X3 clkbuf_leaf_118_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_118_clk));
 CLKBUF_X3 clkbuf_leaf_119_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_119_clk));
 CLKBUF_X3 clkbuf_leaf_120_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_120_clk));
 CLKBUF_X3 clkbuf_leaf_121_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_121_clk));
 CLKBUF_X3 clkbuf_leaf_122_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_122_clk));
 CLKBUF_X3 clkbuf_leaf_123_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_123_clk));
 CLKBUF_X3 clkbuf_leaf_124_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_124_clk));
 CLKBUF_X3 clkbuf_leaf_125_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_125_clk));
 CLKBUF_X3 clkbuf_leaf_126_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_126_clk));
 CLKBUF_X3 clkbuf_leaf_127_clk (.A(clknet_4_7_0_clk),
    .Z(clknet_leaf_127_clk));
 CLKBUF_X3 clkbuf_leaf_128_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_128_clk));
 CLKBUF_X3 clkbuf_leaf_129_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_129_clk));
 CLKBUF_X3 clkbuf_leaf_130_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_130_clk));
 CLKBUF_X3 clkbuf_leaf_131_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_131_clk));
 CLKBUF_X3 clkbuf_leaf_132_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_132_clk));
 CLKBUF_X3 clkbuf_leaf_133_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_133_clk));
 CLKBUF_X3 clkbuf_leaf_134_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_134_clk));
 CLKBUF_X3 clkbuf_leaf_135_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_135_clk));
 CLKBUF_X3 clkbuf_leaf_136_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_136_clk));
 CLKBUF_X3 clkbuf_leaf_137_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_137_clk));
 CLKBUF_X3 clkbuf_leaf_138_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_138_clk));
 CLKBUF_X3 clkbuf_leaf_139_clk (.A(clknet_4_5_0_clk),
    .Z(clknet_leaf_139_clk));
 CLKBUF_X3 clkbuf_leaf_140_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_140_clk));
 CLKBUF_X3 clkbuf_leaf_141_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_141_clk));
 CLKBUF_X3 clkbuf_leaf_142_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_142_clk));
 CLKBUF_X3 clkbuf_leaf_143_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_143_clk));
 CLKBUF_X3 clkbuf_leaf_144_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_144_clk));
 CLKBUF_X3 clkbuf_leaf_145_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_145_clk));
 CLKBUF_X3 clkbuf_leaf_146_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_146_clk));
 CLKBUF_X3 clkbuf_leaf_147_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_147_clk));
 CLKBUF_X3 clkbuf_leaf_148_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_148_clk));
 CLKBUF_X3 clkbuf_leaf_149_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_149_clk));
 CLKBUF_X3 clkbuf_leaf_150_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_150_clk));
 CLKBUF_X3 clkbuf_leaf_151_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_151_clk));
 CLKBUF_X3 clkbuf_leaf_152_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_152_clk));
 CLKBUF_X3 clkbuf_leaf_153_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_153_clk));
 CLKBUF_X3 clkbuf_leaf_154_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_154_clk));
 CLKBUF_X3 clkbuf_leaf_155_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_155_clk));
 CLKBUF_X3 clkbuf_leaf_156_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_156_clk));
 CLKBUF_X3 clkbuf_leaf_157_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_157_clk));
 CLKBUF_X3 clkbuf_leaf_158_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_158_clk));
 CLKBUF_X3 clkbuf_leaf_159_clk (.A(clknet_4_6_0_clk),
    .Z(clknet_leaf_159_clk));
 CLKBUF_X3 clkbuf_leaf_160_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_160_clk));
 CLKBUF_X3 clkbuf_leaf_161_clk (.A(clknet_4_3_0_clk),
    .Z(clknet_leaf_161_clk));
 CLKBUF_X3 clkbuf_leaf_162_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_162_clk));
 CLKBUF_X3 clkbuf_leaf_163_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_163_clk));
 CLKBUF_X3 clkbuf_leaf_164_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_164_clk));
 CLKBUF_X3 clkbuf_leaf_165_clk (.A(clknet_4_4_0_clk),
    .Z(clknet_leaf_165_clk));
 CLKBUF_X3 clkbuf_leaf_166_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_166_clk));
 CLKBUF_X3 clkbuf_leaf_167_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_167_clk));
 CLKBUF_X3 clkbuf_leaf_168_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_168_clk));
 CLKBUF_X3 clkbuf_leaf_169_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_169_clk));
 CLKBUF_X3 clkbuf_leaf_170_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_170_clk));
 CLKBUF_X3 clkbuf_leaf_171_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_171_clk));
 CLKBUF_X3 clkbuf_leaf_172_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_172_clk));
 CLKBUF_X3 clkbuf_leaf_173_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_173_clk));
 CLKBUF_X3 clkbuf_leaf_174_clk (.A(clknet_4_1_0_clk),
    .Z(clknet_leaf_174_clk));
 CLKBUF_X3 clkbuf_leaf_175_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_175_clk));
 CLKBUF_X3 clkbuf_leaf_176_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_176_clk));
 CLKBUF_X3 clkbuf_leaf_177_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_177_clk));
 CLKBUF_X3 clkbuf_leaf_178_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_178_clk));
 CLKBUF_X3 clkbuf_leaf_179_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_179_clk));
 CLKBUF_X3 clkbuf_leaf_180_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_180_clk));
 CLKBUF_X3 clkbuf_leaf_181_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_181_clk));
 CLKBUF_X3 clkbuf_leaf_182_clk (.A(clknet_4_0_0_clk),
    .Z(clknet_leaf_182_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X4 clkload0 (.A(clknet_4_0_0_clk));
 INV_X2 clkload1 (.A(clknet_4_1_0_clk));
 CLKBUF_X3 clkload2 (.A(clknet_4_2_0_clk));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk));
 INV_X4 clkload4 (.A(clknet_4_4_0_clk));
 INV_X2 clkload5 (.A(clknet_4_5_0_clk));
 INV_X2 clkload6 (.A(clknet_4_6_0_clk));
 INV_X4 clkload7 (.A(clknet_4_7_0_clk));
 INV_X2 clkload8 (.A(clknet_4_8_0_clk));
 INV_X4 clkload9 (.A(clknet_4_9_0_clk));
 INV_X2 clkload10 (.A(clknet_4_10_0_clk));
 INV_X4 clkload11 (.A(clknet_4_11_0_clk));
 INV_X4 clkload12 (.A(clknet_4_12_0_clk));
 INV_X4 clkload13 (.A(clknet_4_13_0_clk));
 INV_X2 clkload14 (.A(clknet_4_14_0_clk));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_2_clk));
 INV_X2 clkload16 (.A(clknet_leaf_3_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_175_clk));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_176_clk));
 CLKBUF_X1 clkload19 (.A(clknet_leaf_177_clk));
 INV_X1 clkload20 (.A(clknet_leaf_178_clk));
 INV_X1 clkload21 (.A(clknet_leaf_179_clk));
 INV_X2 clkload22 (.A(clknet_leaf_181_clk));
 INV_X1 clkload23 (.A(clknet_leaf_182_clk));
 INV_X1 clkload24 (.A(clknet_leaf_162_clk));
 INV_X2 clkload25 (.A(clknet_leaf_163_clk));
 INV_X1 clkload26 (.A(clknet_leaf_164_clk));
 INV_X2 clkload27 (.A(clknet_leaf_166_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_167_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_168_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_169_clk));
 INV_X2 clkload31 (.A(clknet_leaf_170_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_171_clk));
 INV_X1 clkload33 (.A(clknet_leaf_172_clk));
 INV_X1 clkload34 (.A(clknet_leaf_174_clk));
 INV_X1 clkload35 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_1_clk));
 INV_X4 clkload37 (.A(clknet_leaf_4_clk));
 INV_X1 clkload38 (.A(clknet_leaf_5_clk));
 INV_X1 clkload39 (.A(clknet_leaf_7_clk));
 INV_X1 clkload40 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload41 (.A(clknet_leaf_9_clk));
 INV_X4 clkload42 (.A(clknet_leaf_10_clk));
 INV_X1 clkload43 (.A(clknet_leaf_11_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_12_clk));
 CLKBUF_X1 clkload45 (.A(clknet_leaf_13_clk));
 INV_X2 clkload46 (.A(clknet_leaf_14_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_18_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_19_clk));
 INV_X2 clkload49 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_21_clk));
 INV_X2 clkload51 (.A(clknet_leaf_22_clk));
 INV_X4 clkload52 (.A(clknet_leaf_160_clk));
 INV_X1 clkload53 (.A(clknet_leaf_161_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_140_clk));
 INV_X1 clkload55 (.A(clknet_leaf_144_clk));
 INV_X1 clkload56 (.A(clknet_leaf_145_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_146_clk));
 INV_X4 clkload58 (.A(clknet_leaf_147_clk));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_148_clk));
 INV_X2 clkload60 (.A(clknet_leaf_149_clk));
 INV_X2 clkload61 (.A(clknet_leaf_165_clk));
 INV_X2 clkload62 (.A(clknet_leaf_128_clk));
 INV_X2 clkload63 (.A(clknet_leaf_129_clk));
 INV_X4 clkload64 (.A(clknet_leaf_130_clk));
 INV_X2 clkload65 (.A(clknet_leaf_131_clk));
 INV_X1 clkload66 (.A(clknet_leaf_132_clk));
 INV_X1 clkload67 (.A(clknet_leaf_133_clk));
 INV_X1 clkload68 (.A(clknet_leaf_134_clk));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_135_clk));
 INV_X2 clkload70 (.A(clknet_leaf_136_clk));
 INV_X1 clkload71 (.A(clknet_leaf_138_clk));
 INV_X2 clkload72 (.A(clknet_leaf_139_clk));
 INV_X1 clkload73 (.A(clknet_leaf_116_clk));
 INV_X2 clkload74 (.A(clknet_leaf_117_clk));
 CLKBUF_X1 clkload75 (.A(clknet_leaf_151_clk));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_152_clk));
 INV_X1 clkload77 (.A(clknet_leaf_153_clk));
 INV_X1 clkload78 (.A(clknet_leaf_155_clk));
 INV_X2 clkload79 (.A(clknet_leaf_157_clk));
 CLKBUF_X1 clkload80 (.A(clknet_leaf_158_clk));
 INV_X1 clkload81 (.A(clknet_leaf_159_clk));
 CLKBUF_X1 clkload82 (.A(clknet_leaf_118_clk));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_119_clk));
 CLKBUF_X1 clkload84 (.A(clknet_leaf_120_clk));
 CLKBUF_X1 clkload85 (.A(clknet_leaf_121_clk));
 INV_X1 clkload86 (.A(clknet_leaf_122_clk));
 CLKBUF_X1 clkload87 (.A(clknet_leaf_123_clk));
 INV_X2 clkload88 (.A(clknet_leaf_124_clk));
 INV_X2 clkload89 (.A(clknet_leaf_126_clk));
 INV_X1 clkload90 (.A(clknet_leaf_127_clk));
 CLKBUF_X1 clkload91 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload92 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload93 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload94 (.A(clknet_leaf_35_clk));
 INV_X2 clkload95 (.A(clknet_leaf_36_clk));
 INV_X2 clkload96 (.A(clknet_leaf_37_clk));
 INV_X2 clkload97 (.A(clknet_leaf_38_clk));
 INV_X1 clkload98 (.A(clknet_leaf_39_clk));
 INV_X1 clkload99 (.A(clknet_leaf_42_clk));
 INV_X1 clkload100 (.A(clknet_leaf_44_clk));
 INV_X1 clkload101 (.A(clknet_leaf_23_clk));
 INV_X1 clkload102 (.A(clknet_leaf_24_clk));
 INV_X2 clkload103 (.A(clknet_leaf_25_clk));
 INV_X2 clkload104 (.A(clknet_leaf_26_clk));
 INV_X2 clkload105 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload106 (.A(clknet_leaf_28_clk));
 INV_X4 clkload107 (.A(clknet_leaf_29_clk));
 INV_X2 clkload108 (.A(clknet_leaf_69_clk));
 INV_X2 clkload109 (.A(clknet_leaf_70_clk));
 INV_X1 clkload110 (.A(clknet_leaf_41_clk));
 INV_X2 clkload111 (.A(clknet_leaf_45_clk));
 INV_X1 clkload112 (.A(clknet_leaf_47_clk));
 INV_X1 clkload113 (.A(clknet_leaf_48_clk));
 INV_X2 clkload114 (.A(clknet_leaf_49_clk));
 INV_X1 clkload115 (.A(clknet_leaf_50_clk));
 INV_X2 clkload116 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload117 (.A(clknet_leaf_52_clk));
 CLKBUF_X1 clkload118 (.A(clknet_leaf_53_clk));
 CLKBUF_X1 clkload119 (.A(clknet_leaf_54_clk));
 INV_X1 clkload120 (.A(clknet_leaf_56_clk));
 INV_X1 clkload121 (.A(clknet_leaf_57_clk));
 INV_X1 clkload122 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload123 (.A(clknet_leaf_60_clk));
 CLKBUF_X1 clkload124 (.A(clknet_leaf_65_clk));
 INV_X1 clkload125 (.A(clknet_leaf_66_clk));
 CLKBUF_X1 clkload126 (.A(clknet_leaf_67_clk));
 INV_X2 clkload127 (.A(clknet_leaf_68_clk));
 CLKBUF_X1 clkload128 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload129 (.A(clknet_leaf_73_clk));
 INV_X2 clkload130 (.A(clknet_leaf_74_clk));
 INV_X2 clkload131 (.A(clknet_leaf_75_clk));
 INV_X2 clkload132 (.A(clknet_leaf_76_clk));
 INV_X2 clkload133 (.A(clknet_leaf_77_clk));
 INV_X1 clkload134 (.A(clknet_leaf_112_clk));
 INV_X2 clkload135 (.A(clknet_leaf_113_clk));
 INV_X2 clkload136 (.A(clknet_leaf_114_clk));
 INV_X2 clkload137 (.A(clknet_leaf_115_clk));
 CLKBUF_X1 clkload138 (.A(clknet_leaf_78_clk));
 CLKBUF_X1 clkload139 (.A(clknet_leaf_102_clk));
 CLKBUF_X1 clkload140 (.A(clknet_leaf_103_clk));
 INV_X2 clkload141 (.A(clknet_leaf_104_clk));
 INV_X2 clkload142 (.A(clknet_leaf_105_clk));
 CLKBUF_X1 clkload143 (.A(clknet_leaf_106_clk));
 CLKBUF_X1 clkload144 (.A(clknet_leaf_109_clk));
 CLKBUF_X1 clkload145 (.A(clknet_leaf_110_clk));
 CLKBUF_X1 clkload146 (.A(clknet_leaf_111_clk));
 INV_X1 clkload147 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload148 (.A(clknet_leaf_62_clk));
 INV_X4 clkload149 (.A(clknet_leaf_63_clk));
 INV_X1 clkload150 (.A(clknet_leaf_82_clk));
 INV_X2 clkload151 (.A(clknet_leaf_84_clk));
 INV_X4 clkload152 (.A(clknet_leaf_85_clk));
 CLKBUF_X1 clkload153 (.A(clknet_leaf_88_clk));
 CLKBUF_X1 clkload154 (.A(clknet_leaf_79_clk));
 CLKBUF_X1 clkload155 (.A(clknet_leaf_89_clk));
 CLKBUF_X1 clkload156 (.A(clknet_leaf_90_clk));
 CLKBUF_X1 clkload157 (.A(clknet_leaf_92_clk));
 INV_X2 clkload158 (.A(clknet_leaf_93_clk));
 CLKBUF_X1 clkload159 (.A(clknet_leaf_95_clk));
 INV_X1 clkload160 (.A(clknet_leaf_97_clk));
 INV_X2 clkload161 (.A(clknet_leaf_98_clk));
 CLKBUF_X1 clkload162 (.A(clknet_leaf_99_clk));
 INV_X2 clkload163 (.A(clknet_leaf_100_clk));
 INV_X1 clkload164 (.A(clknet_leaf_101_clk));
 FILLCELL_X8 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_9 ();
 FILLCELL_X1 FILLER_0_11 ();
 FILLCELL_X32 FILLER_0_15 ();
 FILLCELL_X32 FILLER_0_47 ();
 FILLCELL_X32 FILLER_0_79 ();
 FILLCELL_X32 FILLER_0_111 ();
 FILLCELL_X8 FILLER_0_143 ();
 FILLCELL_X4 FILLER_0_151 ();
 FILLCELL_X2 FILLER_0_155 ();
 FILLCELL_X2 FILLER_0_272 ();
 FILLCELL_X1 FILLER_0_302 ();
 FILLCELL_X2 FILLER_0_376 ();
 FILLCELL_X32 FILLER_0_396 ();
 FILLCELL_X16 FILLER_0_428 ();
 FILLCELL_X8 FILLER_0_444 ();
 FILLCELL_X1 FILLER_0_452 ();
 FILLCELL_X4 FILLER_0_456 ();
 FILLCELL_X2 FILLER_0_460 ();
 FILLCELL_X1 FILLER_0_462 ();
 FILLCELL_X2 FILLER_0_466 ();
 FILLCELL_X1 FILLER_0_468 ();
 FILLCELL_X16 FILLER_0_472 ();
 FILLCELL_X1 FILLER_0_488 ();
 FILLCELL_X32 FILLER_0_492 ();
 FILLCELL_X4 FILLER_0_524 ();
 FILLCELL_X4 FILLER_0_531 ();
 FILLCELL_X1 FILLER_0_535 ();
 FILLCELL_X2 FILLER_0_539 ();
 FILLCELL_X1 FILLER_0_541 ();
 FILLCELL_X4 FILLER_0_548 ();
 FILLCELL_X2 FILLER_0_552 ();
 FILLCELL_X1 FILLER_0_584 ();
 FILLCELL_X4 FILLER_0_599 ();
 FILLCELL_X2 FILLER_0_621 ();
 FILLCELL_X1 FILLER_0_623 ();
 FILLCELL_X4 FILLER_0_627 ();
 FILLCELL_X4 FILLER_0_642 ();
 FILLCELL_X4 FILLER_0_649 ();
 FILLCELL_X4 FILLER_0_659 ();
 FILLCELL_X2 FILLER_0_663 ();
 FILLCELL_X4 FILLER_0_668 ();
 FILLCELL_X2 FILLER_0_672 ();
 FILLCELL_X2 FILLER_0_684 ();
 FILLCELL_X8 FILLER_0_690 ();
 FILLCELL_X2 FILLER_0_698 ();
 FILLCELL_X4 FILLER_0_703 ();
 FILLCELL_X2 FILLER_0_707 ();
 FILLCELL_X4 FILLER_0_713 ();
 FILLCELL_X1 FILLER_0_731 ();
 FILLCELL_X1 FILLER_0_736 ();
 FILLCELL_X1 FILLER_0_744 ();
 FILLCELL_X4 FILLER_0_748 ();
 FILLCELL_X2 FILLER_0_752 ();
 FILLCELL_X1 FILLER_0_754 ();
 FILLCELL_X2 FILLER_0_758 ();
 FILLCELL_X1 FILLER_0_760 ();
 FILLCELL_X4 FILLER_0_765 ();
 FILLCELL_X1 FILLER_0_769 ();
 FILLCELL_X4 FILLER_0_773 ();
 FILLCELL_X2 FILLER_0_777 ();
 FILLCELL_X1 FILLER_0_779 ();
 FILLCELL_X2 FILLER_0_787 ();
 FILLCELL_X2 FILLER_0_793 ();
 FILLCELL_X1 FILLER_0_795 ();
 FILLCELL_X4 FILLER_0_806 ();
 FILLCELL_X2 FILLER_0_810 ();
 FILLCELL_X32 FILLER_0_834 ();
 FILLCELL_X32 FILLER_0_866 ();
 FILLCELL_X2 FILLER_0_898 ();
 FILLCELL_X4 FILLER_0_932 ();
 FILLCELL_X2 FILLER_0_965 ();
 FILLCELL_X2 FILLER_0_1007 ();
 FILLCELL_X1 FILLER_0_1009 ();
 FILLCELL_X8 FILLER_0_1032 ();
 FILLCELL_X4 FILLER_0_1040 ();
 FILLCELL_X2 FILLER_0_1044 ();
 FILLCELL_X1 FILLER_0_1046 ();
 FILLCELL_X1 FILLER_0_1050 ();
 FILLCELL_X1 FILLER_0_1054 ();
 FILLCELL_X2 FILLER_0_1059 ();
 FILLCELL_X16 FILLER_0_1127 ();
 FILLCELL_X4 FILLER_0_1143 ();
 FILLCELL_X1 FILLER_0_1147 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X8 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_157 ();
 FILLCELL_X2 FILLER_1_190 ();
 FILLCELL_X32 FILLER_1_195 ();
 FILLCELL_X8 FILLER_1_227 ();
 FILLCELL_X4 FILLER_1_235 ();
 FILLCELL_X2 FILLER_1_239 ();
 FILLCELL_X2 FILLER_1_259 ();
 FILLCELL_X2 FILLER_1_268 ();
 FILLCELL_X4 FILLER_1_391 ();
 FILLCELL_X1 FILLER_1_395 ();
 FILLCELL_X4 FILLER_1_402 ();
 FILLCELL_X2 FILLER_1_406 ();
 FILLCELL_X32 FILLER_1_430 ();
 FILLCELL_X8 FILLER_1_462 ();
 FILLCELL_X1 FILLER_1_470 ();
 FILLCELL_X32 FILLER_1_477 ();
 FILLCELL_X32 FILLER_1_509 ();
 FILLCELL_X16 FILLER_1_541 ();
 FILLCELL_X4 FILLER_1_557 ();
 FILLCELL_X2 FILLER_1_561 ();
 FILLCELL_X1 FILLER_1_563 ();
 FILLCELL_X1 FILLER_1_609 ();
 FILLCELL_X1 FILLER_1_618 ();
 FILLCELL_X4 FILLER_1_650 ();
 FILLCELL_X8 FILLER_1_658 ();
 FILLCELL_X2 FILLER_1_666 ();
 FILLCELL_X1 FILLER_1_668 ();
 FILLCELL_X4 FILLER_1_674 ();
 FILLCELL_X2 FILLER_1_678 ();
 FILLCELL_X4 FILLER_1_684 ();
 FILLCELL_X2 FILLER_1_688 ();
 FILLCELL_X1 FILLER_1_690 ();
 FILLCELL_X2 FILLER_1_733 ();
 FILLCELL_X16 FILLER_1_755 ();
 FILLCELL_X8 FILLER_1_771 ();
 FILLCELL_X1 FILLER_1_779 ();
 FILLCELL_X8 FILLER_1_800 ();
 FILLCELL_X4 FILLER_1_808 ();
 FILLCELL_X32 FILLER_1_850 ();
 FILLCELL_X16 FILLER_1_882 ();
 FILLCELL_X8 FILLER_1_898 ();
 FILLCELL_X4 FILLER_1_906 ();
 FILLCELL_X1 FILLER_1_910 ();
 FILLCELL_X4 FILLER_1_992 ();
 FILLCELL_X1 FILLER_1_1004 ();
 FILLCELL_X1 FILLER_1_1009 ();
 FILLCELL_X2 FILLER_1_1013 ();
 FILLCELL_X1 FILLER_1_1058 ();
 FILLCELL_X16 FILLER_1_1124 ();
 FILLCELL_X8 FILLER_1_1140 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_81 ();
 FILLCELL_X4 FILLER_2_89 ();
 FILLCELL_X2 FILLER_2_93 ();
 FILLCELL_X1 FILLER_2_95 ();
 FILLCELL_X4 FILLER_2_112 ();
 FILLCELL_X8 FILLER_2_140 ();
 FILLCELL_X4 FILLER_2_148 ();
 FILLCELL_X2 FILLER_2_152 ();
 FILLCELL_X1 FILLER_2_156 ();
 FILLCELL_X2 FILLER_2_185 ();
 FILLCELL_X1 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_287 ();
 FILLCELL_X1 FILLER_2_341 ();
 FILLCELL_X32 FILLER_2_420 ();
 FILLCELL_X32 FILLER_2_452 ();
 FILLCELL_X32 FILLER_2_504 ();
 FILLCELL_X16 FILLER_2_536 ();
 FILLCELL_X4 FILLER_2_552 ();
 FILLCELL_X1 FILLER_2_556 ();
 FILLCELL_X1 FILLER_2_585 ();
 FILLCELL_X1 FILLER_2_588 ();
 FILLCELL_X1 FILLER_2_592 ();
 FILLCELL_X1 FILLER_2_599 ();
 FILLCELL_X2 FILLER_2_604 ();
 FILLCELL_X1 FILLER_2_626 ();
 FILLCELL_X1 FILLER_2_639 ();
 FILLCELL_X8 FILLER_2_658 ();
 FILLCELL_X2 FILLER_2_666 ();
 FILLCELL_X8 FILLER_2_672 ();
 FILLCELL_X2 FILLER_2_680 ();
 FILLCELL_X2 FILLER_2_686 ();
 FILLCELL_X1 FILLER_2_688 ();
 FILLCELL_X2 FILLER_2_693 ();
 FILLCELL_X1 FILLER_2_695 ();
 FILLCELL_X2 FILLER_2_698 ();
 FILLCELL_X1 FILLER_2_709 ();
 FILLCELL_X8 FILLER_2_726 ();
 FILLCELL_X1 FILLER_2_734 ();
 FILLCELL_X4 FILLER_2_769 ();
 FILLCELL_X2 FILLER_2_773 ();
 FILLCELL_X4 FILLER_2_779 ();
 FILLCELL_X2 FILLER_2_783 ();
 FILLCELL_X4 FILLER_2_791 ();
 FILLCELL_X2 FILLER_2_795 ();
 FILLCELL_X1 FILLER_2_813 ();
 FILLCELL_X16 FILLER_2_822 ();
 FILLCELL_X2 FILLER_2_838 ();
 FILLCELL_X16 FILLER_2_872 ();
 FILLCELL_X4 FILLER_2_888 ();
 FILLCELL_X1 FILLER_2_892 ();
 FILLCELL_X1 FILLER_2_913 ();
 FILLCELL_X1 FILLER_2_922 ();
 FILLCELL_X4 FILLER_2_926 ();
 FILLCELL_X2 FILLER_2_930 ();
 FILLCELL_X1 FILLER_2_932 ();
 FILLCELL_X4 FILLER_2_945 ();
 FILLCELL_X1 FILLER_2_949 ();
 FILLCELL_X1 FILLER_2_977 ();
 FILLCELL_X4 FILLER_2_987 ();
 FILLCELL_X1 FILLER_2_991 ();
 FILLCELL_X1 FILLER_2_996 ();
 FILLCELL_X2 FILLER_2_1017 ();
 FILLCELL_X2 FILLER_2_1032 ();
 FILLCELL_X2 FILLER_2_1038 ();
 FILLCELL_X2 FILLER_2_1079 ();
 FILLCELL_X2 FILLER_2_1098 ();
 FILLCELL_X1 FILLER_2_1103 ();
 FILLCELL_X4 FILLER_2_1115 ();
 FILLCELL_X8 FILLER_2_1133 ();
 FILLCELL_X4 FILLER_2_1141 ();
 FILLCELL_X2 FILLER_2_1145 ();
 FILLCELL_X1 FILLER_2_1147 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_97 ();
 FILLCELL_X2 FILLER_3_101 ();
 FILLCELL_X1 FILLER_3_103 ();
 FILLCELL_X16 FILLER_3_106 ();
 FILLCELL_X1 FILLER_3_122 ();
 FILLCELL_X1 FILLER_3_155 ();
 FILLCELL_X1 FILLER_3_158 ();
 FILLCELL_X1 FILLER_3_175 ();
 FILLCELL_X1 FILLER_3_192 ();
 FILLCELL_X2 FILLER_3_248 ();
 FILLCELL_X1 FILLER_3_250 ();
 FILLCELL_X1 FILLER_3_277 ();
 FILLCELL_X2 FILLER_3_290 ();
 FILLCELL_X2 FILLER_3_365 ();
 FILLCELL_X4 FILLER_3_413 ();
 FILLCELL_X16 FILLER_3_439 ();
 FILLCELL_X4 FILLER_3_455 ();
 FILLCELL_X2 FILLER_3_459 ();
 FILLCELL_X1 FILLER_3_461 ();
 FILLCELL_X16 FILLER_3_468 ();
 FILLCELL_X2 FILLER_3_484 ();
 FILLCELL_X4 FILLER_3_492 ();
 FILLCELL_X32 FILLER_3_499 ();
 FILLCELL_X32 FILLER_3_531 ();
 FILLCELL_X2 FILLER_3_619 ();
 FILLCELL_X4 FILLER_3_628 ();
 FILLCELL_X2 FILLER_3_632 ();
 FILLCELL_X1 FILLER_3_634 ();
 FILLCELL_X4 FILLER_3_643 ();
 FILLCELL_X2 FILLER_3_647 ();
 FILLCELL_X1 FILLER_3_649 ();
 FILLCELL_X8 FILLER_3_654 ();
 FILLCELL_X1 FILLER_3_662 ();
 FILLCELL_X4 FILLER_3_667 ();
 FILLCELL_X2 FILLER_3_671 ();
 FILLCELL_X1 FILLER_3_673 ();
 FILLCELL_X2 FILLER_3_678 ();
 FILLCELL_X1 FILLER_3_680 ();
 FILLCELL_X2 FILLER_3_723 ();
 FILLCELL_X2 FILLER_3_771 ();
 FILLCELL_X2 FILLER_3_795 ();
 FILLCELL_X2 FILLER_3_804 ();
 FILLCELL_X1 FILLER_3_806 ();
 FILLCELL_X8 FILLER_3_893 ();
 FILLCELL_X2 FILLER_3_901 ();
 FILLCELL_X2 FILLER_3_946 ();
 FILLCELL_X2 FILLER_3_968 ();
 FILLCELL_X1 FILLER_3_1020 ();
 FILLCELL_X16 FILLER_3_1132 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X2 FILLER_4_49 ();
 FILLCELL_X32 FILLER_4_54 ();
 FILLCELL_X16 FILLER_4_86 ();
 FILLCELL_X4 FILLER_4_102 ();
 FILLCELL_X1 FILLER_4_106 ();
 FILLCELL_X2 FILLER_4_127 ();
 FILLCELL_X1 FILLER_4_147 ();
 FILLCELL_X1 FILLER_4_221 ();
 FILLCELL_X2 FILLER_4_226 ();
 FILLCELL_X1 FILLER_4_260 ();
 FILLCELL_X1 FILLER_4_283 ();
 FILLCELL_X1 FILLER_4_373 ();
 FILLCELL_X1 FILLER_4_380 ();
 FILLCELL_X1 FILLER_4_397 ();
 FILLCELL_X32 FILLER_4_418 ();
 FILLCELL_X32 FILLER_4_452 ();
 FILLCELL_X32 FILLER_4_507 ();
 FILLCELL_X8 FILLER_4_539 ();
 FILLCELL_X4 FILLER_4_547 ();
 FILLCELL_X2 FILLER_4_551 ();
 FILLCELL_X1 FILLER_4_553 ();
 FILLCELL_X8 FILLER_4_556 ();
 FILLCELL_X2 FILLER_4_564 ();
 FILLCELL_X2 FILLER_4_568 ();
 FILLCELL_X4 FILLER_4_572 ();
 FILLCELL_X1 FILLER_4_576 ();
 FILLCELL_X2 FILLER_4_591 ();
 FILLCELL_X4 FILLER_4_595 ();
 FILLCELL_X4 FILLER_4_648 ();
 FILLCELL_X16 FILLER_4_658 ();
 FILLCELL_X2 FILLER_4_674 ();
 FILLCELL_X1 FILLER_4_676 ();
 FILLCELL_X1 FILLER_4_693 ();
 FILLCELL_X8 FILLER_4_698 ();
 FILLCELL_X1 FILLER_4_706 ();
 FILLCELL_X8 FILLER_4_752 ();
 FILLCELL_X1 FILLER_4_760 ();
 FILLCELL_X1 FILLER_4_779 ();
 FILLCELL_X4 FILLER_4_784 ();
 FILLCELL_X1 FILLER_4_788 ();
 FILLCELL_X1 FILLER_4_827 ();
 FILLCELL_X4 FILLER_4_850 ();
 FILLCELL_X1 FILLER_4_854 ();
 FILLCELL_X4 FILLER_4_857 ();
 FILLCELL_X2 FILLER_4_887 ();
 FILLCELL_X16 FILLER_4_893 ();
 FILLCELL_X4 FILLER_4_909 ();
 FILLCELL_X1 FILLER_4_913 ();
 FILLCELL_X2 FILLER_4_916 ();
 FILLCELL_X1 FILLER_4_918 ();
 FILLCELL_X16 FILLER_4_942 ();
 FILLCELL_X4 FILLER_4_958 ();
 FILLCELL_X1 FILLER_4_962 ();
 FILLCELL_X4 FILLER_4_967 ();
 FILLCELL_X2 FILLER_4_986 ();
 FILLCELL_X1 FILLER_4_988 ();
 FILLCELL_X1 FILLER_4_992 ();
 FILLCELL_X2 FILLER_4_1013 ();
 FILLCELL_X1 FILLER_4_1015 ();
 FILLCELL_X1 FILLER_4_1046 ();
 FILLCELL_X2 FILLER_4_1124 ();
 FILLCELL_X1 FILLER_4_1126 ();
 FILLCELL_X16 FILLER_4_1132 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_73 ();
 FILLCELL_X2 FILLER_5_77 ();
 FILLCELL_X1 FILLER_5_103 ();
 FILLCELL_X16 FILLER_5_110 ();
 FILLCELL_X8 FILLER_5_160 ();
 FILLCELL_X2 FILLER_5_168 ();
 FILLCELL_X1 FILLER_5_170 ();
 FILLCELL_X2 FILLER_5_173 ();
 FILLCELL_X1 FILLER_5_175 ();
 FILLCELL_X4 FILLER_5_178 ();
 FILLCELL_X4 FILLER_5_202 ();
 FILLCELL_X1 FILLER_5_206 ();
 FILLCELL_X2 FILLER_5_209 ();
 FILLCELL_X1 FILLER_5_231 ();
 FILLCELL_X1 FILLER_5_262 ();
 FILLCELL_X1 FILLER_5_298 ();
 FILLCELL_X1 FILLER_5_327 ();
 FILLCELL_X4 FILLER_5_352 ();
 FILLCELL_X1 FILLER_5_376 ();
 FILLCELL_X1 FILLER_5_411 ();
 FILLCELL_X1 FILLER_5_434 ();
 FILLCELL_X1 FILLER_5_454 ();
 FILLCELL_X2 FILLER_5_459 ();
 FILLCELL_X1 FILLER_5_461 ();
 FILLCELL_X2 FILLER_5_467 ();
 FILLCELL_X1 FILLER_5_475 ();
 FILLCELL_X2 FILLER_5_501 ();
 FILLCELL_X16 FILLER_5_525 ();
 FILLCELL_X4 FILLER_5_541 ();
 FILLCELL_X1 FILLER_5_545 ();
 FILLCELL_X1 FILLER_5_602 ();
 FILLCELL_X1 FILLER_5_607 ();
 FILLCELL_X1 FILLER_5_612 ();
 FILLCELL_X1 FILLER_5_629 ();
 FILLCELL_X1 FILLER_5_658 ();
 FILLCELL_X4 FILLER_5_661 ();
 FILLCELL_X2 FILLER_5_665 ();
 FILLCELL_X1 FILLER_5_667 ();
 FILLCELL_X4 FILLER_5_720 ();
 FILLCELL_X1 FILLER_5_724 ();
 FILLCELL_X2 FILLER_5_729 ();
 FILLCELL_X1 FILLER_5_731 ();
 FILLCELL_X4 FILLER_5_736 ();
 FILLCELL_X4 FILLER_5_742 ();
 FILLCELL_X4 FILLER_5_748 ();
 FILLCELL_X1 FILLER_5_756 ();
 FILLCELL_X1 FILLER_5_759 ();
 FILLCELL_X1 FILLER_5_770 ();
 FILLCELL_X1 FILLER_5_778 ();
 FILLCELL_X8 FILLER_5_802 ();
 FILLCELL_X2 FILLER_5_810 ();
 FILLCELL_X1 FILLER_5_815 ();
 FILLCELL_X2 FILLER_5_818 ();
 FILLCELL_X1 FILLER_5_824 ();
 FILLCELL_X1 FILLER_5_835 ();
 FILLCELL_X4 FILLER_5_865 ();
 FILLCELL_X2 FILLER_5_869 ();
 FILLCELL_X16 FILLER_5_895 ();
 FILLCELL_X4 FILLER_5_911 ();
 FILLCELL_X1 FILLER_5_915 ();
 FILLCELL_X16 FILLER_5_939 ();
 FILLCELL_X8 FILLER_5_955 ();
 FILLCELL_X4 FILLER_5_963 ();
 FILLCELL_X1 FILLER_5_967 ();
 FILLCELL_X1 FILLER_5_976 ();
 FILLCELL_X1 FILLER_5_981 ();
 FILLCELL_X1 FILLER_5_991 ();
 FILLCELL_X1 FILLER_5_1012 ();
 FILLCELL_X1 FILLER_5_1097 ();
 FILLCELL_X1 FILLER_5_1127 ();
 FILLCELL_X2 FILLER_5_1131 ();
 FILLCELL_X8 FILLER_5_1138 ();
 FILLCELL_X2 FILLER_5_1146 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X2 FILLER_6_65 ();
 FILLCELL_X1 FILLER_6_67 ();
 FILLCELL_X2 FILLER_6_70 ();
 FILLCELL_X1 FILLER_6_88 ();
 FILLCELL_X1 FILLER_6_105 ();
 FILLCELL_X1 FILLER_6_108 ();
 FILLCELL_X1 FILLER_6_141 ();
 FILLCELL_X1 FILLER_6_172 ();
 FILLCELL_X2 FILLER_6_215 ();
 FILLCELL_X4 FILLER_6_219 ();
 FILLCELL_X2 FILLER_6_223 ();
 FILLCELL_X1 FILLER_6_227 ();
 FILLCELL_X1 FILLER_6_232 ();
 FILLCELL_X1 FILLER_6_241 ();
 FILLCELL_X4 FILLER_6_303 ();
 FILLCELL_X1 FILLER_6_307 ();
 FILLCELL_X2 FILLER_6_311 ();
 FILLCELL_X8 FILLER_6_335 ();
 FILLCELL_X1 FILLER_6_376 ();
 FILLCELL_X2 FILLER_6_416 ();
 FILLCELL_X1 FILLER_6_418 ();
 FILLCELL_X2 FILLER_6_482 ();
 FILLCELL_X2 FILLER_6_510 ();
 FILLCELL_X16 FILLER_6_515 ();
 FILLCELL_X8 FILLER_6_531 ();
 FILLCELL_X1 FILLER_6_539 ();
 FILLCELL_X1 FILLER_6_556 ();
 FILLCELL_X2 FILLER_6_573 ();
 FILLCELL_X4 FILLER_6_577 ();
 FILLCELL_X4 FILLER_6_585 ();
 FILLCELL_X2 FILLER_6_589 ();
 FILLCELL_X1 FILLER_6_591 ();
 FILLCELL_X1 FILLER_6_613 ();
 FILLCELL_X2 FILLER_6_618 ();
 FILLCELL_X1 FILLER_6_626 ();
 FILLCELL_X1 FILLER_6_630 ();
 FILLCELL_X8 FILLER_6_632 ();
 FILLCELL_X4 FILLER_6_640 ();
 FILLCELL_X2 FILLER_6_644 ();
 FILLCELL_X4 FILLER_6_667 ();
 FILLCELL_X1 FILLER_6_671 ();
 FILLCELL_X2 FILLER_6_688 ();
 FILLCELL_X2 FILLER_6_693 ();
 FILLCELL_X4 FILLER_6_699 ();
 FILLCELL_X1 FILLER_6_703 ();
 FILLCELL_X1 FILLER_6_724 ();
 FILLCELL_X2 FILLER_6_789 ();
 FILLCELL_X2 FILLER_6_793 ();
 FILLCELL_X1 FILLER_6_795 ();
 FILLCELL_X1 FILLER_6_800 ();
 FILLCELL_X2 FILLER_6_817 ();
 FILLCELL_X1 FILLER_6_823 ();
 FILLCELL_X2 FILLER_6_828 ();
 FILLCELL_X4 FILLER_6_832 ();
 FILLCELL_X1 FILLER_6_840 ();
 FILLCELL_X1 FILLER_6_845 ();
 FILLCELL_X1 FILLER_6_856 ();
 FILLCELL_X1 FILLER_6_873 ();
 FILLCELL_X16 FILLER_6_894 ();
 FILLCELL_X8 FILLER_6_910 ();
 FILLCELL_X4 FILLER_6_918 ();
 FILLCELL_X2 FILLER_6_922 ();
 FILLCELL_X1 FILLER_6_924 ();
 FILLCELL_X16 FILLER_6_945 ();
 FILLCELL_X4 FILLER_6_961 ();
 FILLCELL_X8 FILLER_6_975 ();
 FILLCELL_X4 FILLER_6_983 ();
 FILLCELL_X2 FILLER_6_987 ();
 FILLCELL_X1 FILLER_6_989 ();
 FILLCELL_X4 FILLER_6_1020 ();
 FILLCELL_X4 FILLER_6_1027 ();
 FILLCELL_X2 FILLER_6_1031 ();
 FILLCELL_X1 FILLER_6_1033 ();
 FILLCELL_X1 FILLER_6_1088 ();
 FILLCELL_X1 FILLER_6_1094 ();
 FILLCELL_X1 FILLER_6_1128 ();
 FILLCELL_X16 FILLER_6_1132 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X16 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_49 ();
 FILLCELL_X4 FILLER_7_57 ();
 FILLCELL_X2 FILLER_7_61 ();
 FILLCELL_X2 FILLER_7_137 ();
 FILLCELL_X2 FILLER_7_143 ();
 FILLCELL_X2 FILLER_7_151 ();
 FILLCELL_X1 FILLER_7_157 ();
 FILLCELL_X1 FILLER_7_162 ();
 FILLCELL_X8 FILLER_7_195 ();
 FILLCELL_X2 FILLER_7_203 ();
 FILLCELL_X2 FILLER_7_237 ();
 FILLCELL_X1 FILLER_7_239 ();
 FILLCELL_X2 FILLER_7_256 ();
 FILLCELL_X4 FILLER_7_283 ();
 FILLCELL_X1 FILLER_7_287 ();
 FILLCELL_X2 FILLER_7_291 ();
 FILLCELL_X1 FILLER_7_293 ();
 FILLCELL_X8 FILLER_7_308 ();
 FILLCELL_X4 FILLER_7_320 ();
 FILLCELL_X1 FILLER_7_324 ();
 FILLCELL_X2 FILLER_7_361 ();
 FILLCELL_X1 FILLER_7_380 ();
 FILLCELL_X2 FILLER_7_384 ();
 FILLCELL_X1 FILLER_7_386 ();
 FILLCELL_X1 FILLER_7_413 ();
 FILLCELL_X1 FILLER_7_431 ();
 FILLCELL_X1 FILLER_7_494 ();
 FILLCELL_X16 FILLER_7_527 ();
 FILLCELL_X2 FILLER_7_543 ();
 FILLCELL_X1 FILLER_7_545 ();
 FILLCELL_X1 FILLER_7_578 ();
 FILLCELL_X2 FILLER_7_597 ();
 FILLCELL_X1 FILLER_7_599 ();
 FILLCELL_X1 FILLER_7_603 ();
 FILLCELL_X1 FILLER_7_608 ();
 FILLCELL_X1 FILLER_7_613 ();
 FILLCELL_X1 FILLER_7_634 ();
 FILLCELL_X1 FILLER_7_653 ();
 FILLCELL_X8 FILLER_7_657 ();
 FILLCELL_X4 FILLER_7_665 ();
 FILLCELL_X1 FILLER_7_673 ();
 FILLCELL_X1 FILLER_7_676 ();
 FILLCELL_X2 FILLER_7_685 ();
 FILLCELL_X1 FILLER_7_687 ();
 FILLCELL_X2 FILLER_7_690 ();
 FILLCELL_X8 FILLER_7_701 ();
 FILLCELL_X1 FILLER_7_711 ();
 FILLCELL_X8 FILLER_7_720 ();
 FILLCELL_X4 FILLER_7_736 ();
 FILLCELL_X2 FILLER_7_740 ();
 FILLCELL_X1 FILLER_7_742 ();
 FILLCELL_X1 FILLER_7_750 ();
 FILLCELL_X1 FILLER_7_757 ();
 FILLCELL_X1 FILLER_7_788 ();
 FILLCELL_X1 FILLER_7_793 ();
 FILLCELL_X4 FILLER_7_834 ();
 FILLCELL_X1 FILLER_7_886 ();
 FILLCELL_X32 FILLER_7_901 ();
 FILLCELL_X2 FILLER_7_933 ();
 FILLCELL_X1 FILLER_7_949 ();
 FILLCELL_X1 FILLER_7_957 ();
 FILLCELL_X1 FILLER_7_962 ();
 FILLCELL_X1 FILLER_7_967 ();
 FILLCELL_X4 FILLER_7_982 ();
 FILLCELL_X2 FILLER_7_986 ();
 FILLCELL_X1 FILLER_7_1006 ();
 FILLCELL_X4 FILLER_7_1030 ();
 FILLCELL_X2 FILLER_7_1034 ();
 FILLCELL_X1 FILLER_7_1046 ();
 FILLCELL_X1 FILLER_7_1093 ();
 FILLCELL_X2 FILLER_7_1103 ();
 FILLCELL_X1 FILLER_7_1105 ();
 FILLCELL_X1 FILLER_7_1113 ();
 FILLCELL_X1 FILLER_7_1121 ();
 FILLCELL_X1 FILLER_7_1127 ();
 FILLCELL_X8 FILLER_7_1135 ();
 FILLCELL_X4 FILLER_7_1143 ();
 FILLCELL_X1 FILLER_7_1147 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_9 ();
 FILLCELL_X1 FILLER_8_11 ();
 FILLCELL_X32 FILLER_8_19 ();
 FILLCELL_X16 FILLER_8_51 ();
 FILLCELL_X2 FILLER_8_67 ();
 FILLCELL_X1 FILLER_8_69 ();
 FILLCELL_X1 FILLER_8_95 ();
 FILLCELL_X1 FILLER_8_106 ();
 FILLCELL_X1 FILLER_8_139 ();
 FILLCELL_X4 FILLER_8_160 ();
 FILLCELL_X1 FILLER_8_164 ();
 FILLCELL_X2 FILLER_8_202 ();
 FILLCELL_X2 FILLER_8_207 ();
 FILLCELL_X1 FILLER_8_209 ();
 FILLCELL_X2 FILLER_8_212 ();
 FILLCELL_X1 FILLER_8_220 ();
 FILLCELL_X2 FILLER_8_235 ();
 FILLCELL_X1 FILLER_8_237 ();
 FILLCELL_X2 FILLER_8_258 ();
 FILLCELL_X1 FILLER_8_260 ();
 FILLCELL_X16 FILLER_8_269 ();
 FILLCELL_X8 FILLER_8_285 ();
 FILLCELL_X4 FILLER_8_293 ();
 FILLCELL_X2 FILLER_8_297 ();
 FILLCELL_X2 FILLER_8_329 ();
 FILLCELL_X1 FILLER_8_331 ();
 FILLCELL_X1 FILLER_8_371 ();
 FILLCELL_X1 FILLER_8_418 ();
 FILLCELL_X1 FILLER_8_467 ();
 FILLCELL_X2 FILLER_8_471 ();
 FILLCELL_X1 FILLER_8_494 ();
 FILLCELL_X2 FILLER_8_521 ();
 FILLCELL_X2 FILLER_8_528 ();
 FILLCELL_X4 FILLER_8_535 ();
 FILLCELL_X8 FILLER_8_541 ();
 FILLCELL_X2 FILLER_8_549 ();
 FILLCELL_X1 FILLER_8_551 ();
 FILLCELL_X1 FILLER_8_568 ();
 FILLCELL_X4 FILLER_8_571 ();
 FILLCELL_X2 FILLER_8_575 ();
 FILLCELL_X4 FILLER_8_579 ();
 FILLCELL_X1 FILLER_8_583 ();
 FILLCELL_X4 FILLER_8_626 ();
 FILLCELL_X1 FILLER_8_630 ();
 FILLCELL_X1 FILLER_8_662 ();
 FILLCELL_X2 FILLER_8_681 ();
 FILLCELL_X1 FILLER_8_683 ();
 FILLCELL_X1 FILLER_8_686 ();
 FILLCELL_X8 FILLER_8_755 ();
 FILLCELL_X2 FILLER_8_763 ();
 FILLCELL_X1 FILLER_8_765 ();
 FILLCELL_X1 FILLER_8_804 ();
 FILLCELL_X8 FILLER_8_847 ();
 FILLCELL_X1 FILLER_8_855 ();
 FILLCELL_X2 FILLER_8_883 ();
 FILLCELL_X16 FILLER_8_905 ();
 FILLCELL_X4 FILLER_8_921 ();
 FILLCELL_X2 FILLER_8_925 ();
 FILLCELL_X1 FILLER_8_955 ();
 FILLCELL_X2 FILLER_8_966 ();
 FILLCELL_X1 FILLER_8_968 ();
 FILLCELL_X2 FILLER_8_984 ();
 FILLCELL_X2 FILLER_8_993 ();
 FILLCELL_X1 FILLER_8_995 ();
 FILLCELL_X4 FILLER_8_1008 ();
 FILLCELL_X2 FILLER_8_1012 ();
 FILLCELL_X1 FILLER_8_1014 ();
 FILLCELL_X1 FILLER_8_1035 ();
 FILLCELL_X2 FILLER_8_1048 ();
 FILLCELL_X1 FILLER_8_1068 ();
 FILLCELL_X1 FILLER_8_1080 ();
 FILLCELL_X4 FILLER_8_1142 ();
 FILLCELL_X2 FILLER_8_1146 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X8 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_57 ();
 FILLCELL_X1 FILLER_9_61 ();
 FILLCELL_X1 FILLER_9_109 ();
 FILLCELL_X1 FILLER_9_114 ();
 FILLCELL_X1 FILLER_9_119 ();
 FILLCELL_X1 FILLER_9_124 ();
 FILLCELL_X4 FILLER_9_133 ();
 FILLCELL_X1 FILLER_9_137 ();
 FILLCELL_X4 FILLER_9_140 ();
 FILLCELL_X2 FILLER_9_155 ();
 FILLCELL_X1 FILLER_9_171 ();
 FILLCELL_X2 FILLER_9_224 ();
 FILLCELL_X1 FILLER_9_226 ();
 FILLCELL_X1 FILLER_9_231 ();
 FILLCELL_X2 FILLER_9_239 ();
 FILLCELL_X1 FILLER_9_241 ();
 FILLCELL_X4 FILLER_9_323 ();
 FILLCELL_X2 FILLER_9_327 ();
 FILLCELL_X1 FILLER_9_512 ();
 FILLCELL_X1 FILLER_9_530 ();
 FILLCELL_X16 FILLER_9_543 ();
 FILLCELL_X4 FILLER_9_559 ();
 FILLCELL_X2 FILLER_9_563 ();
 FILLCELL_X4 FILLER_9_581 ();
 FILLCELL_X2 FILLER_9_585 ();
 FILLCELL_X4 FILLER_9_589 ();
 FILLCELL_X4 FILLER_9_597 ();
 FILLCELL_X2 FILLER_9_601 ();
 FILLCELL_X2 FILLER_9_607 ();
 FILLCELL_X1 FILLER_9_612 ();
 FILLCELL_X1 FILLER_9_617 ();
 FILLCELL_X2 FILLER_9_634 ();
 FILLCELL_X2 FILLER_9_638 ();
 FILLCELL_X1 FILLER_9_640 ();
 FILLCELL_X2 FILLER_9_650 ();
 FILLCELL_X1 FILLER_9_668 ();
 FILLCELL_X2 FILLER_9_707 ();
 FILLCELL_X4 FILLER_9_733 ();
 FILLCELL_X2 FILLER_9_737 ();
 FILLCELL_X1 FILLER_9_741 ();
 FILLCELL_X1 FILLER_9_744 ();
 FILLCELL_X2 FILLER_9_749 ();
 FILLCELL_X1 FILLER_9_755 ();
 FILLCELL_X1 FILLER_9_775 ();
 FILLCELL_X4 FILLER_9_778 ();
 FILLCELL_X2 FILLER_9_782 ();
 FILLCELL_X1 FILLER_9_784 ();
 FILLCELL_X4 FILLER_9_803 ();
 FILLCELL_X8 FILLER_9_809 ();
 FILLCELL_X4 FILLER_9_817 ();
 FILLCELL_X4 FILLER_9_901 ();
 FILLCELL_X2 FILLER_9_905 ();
 FILLCELL_X1 FILLER_9_951 ();
 FILLCELL_X4 FILLER_9_982 ();
 FILLCELL_X1 FILLER_9_992 ();
 FILLCELL_X1 FILLER_9_1000 ();
 FILLCELL_X2 FILLER_9_1016 ();
 FILLCELL_X1 FILLER_9_1028 ();
 FILLCELL_X2 FILLER_9_1032 ();
 FILLCELL_X1 FILLER_9_1034 ();
 FILLCELL_X1 FILLER_9_1045 ();
 FILLCELL_X1 FILLER_9_1051 ();
 FILLCELL_X4 FILLER_9_1059 ();
 FILLCELL_X2 FILLER_9_1079 ();
 FILLCELL_X1 FILLER_9_1136 ();
 FILLCELL_X8 FILLER_9_1140 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X16 FILLER_10_33 ();
 FILLCELL_X1 FILLER_10_49 ();
 FILLCELL_X4 FILLER_10_52 ();
 FILLCELL_X4 FILLER_10_74 ();
 FILLCELL_X1 FILLER_10_96 ();
 FILLCELL_X1 FILLER_10_102 ();
 FILLCELL_X8 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_151 ();
 FILLCELL_X1 FILLER_10_155 ();
 FILLCELL_X4 FILLER_10_160 ();
 FILLCELL_X4 FILLER_10_187 ();
 FILLCELL_X2 FILLER_10_191 ();
 FILLCELL_X2 FILLER_10_197 ();
 FILLCELL_X2 FILLER_10_219 ();
 FILLCELL_X1 FILLER_10_225 ();
 FILLCELL_X2 FILLER_10_235 ();
 FILLCELL_X2 FILLER_10_260 ();
 FILLCELL_X2 FILLER_10_292 ();
 FILLCELL_X4 FILLER_10_321 ();
 FILLCELL_X2 FILLER_10_325 ();
 FILLCELL_X1 FILLER_10_327 ();
 FILLCELL_X1 FILLER_10_385 ();
 FILLCELL_X1 FILLER_10_406 ();
 FILLCELL_X1 FILLER_10_448 ();
 FILLCELL_X2 FILLER_10_507 ();
 FILLCELL_X4 FILLER_10_544 ();
 FILLCELL_X2 FILLER_10_548 ();
 FILLCELL_X1 FILLER_10_550 ();
 FILLCELL_X2 FILLER_10_555 ();
 FILLCELL_X1 FILLER_10_557 ();
 FILLCELL_X2 FILLER_10_622 ();
 FILLCELL_X1 FILLER_10_624 ();
 FILLCELL_X2 FILLER_10_628 ();
 FILLCELL_X1 FILLER_10_630 ();
 FILLCELL_X4 FILLER_10_672 ();
 FILLCELL_X1 FILLER_10_676 ();
 FILLCELL_X4 FILLER_10_681 ();
 FILLCELL_X2 FILLER_10_685 ();
 FILLCELL_X1 FILLER_10_703 ();
 FILLCELL_X8 FILLER_10_720 ();
 FILLCELL_X2 FILLER_10_731 ();
 FILLCELL_X2 FILLER_10_768 ();
 FILLCELL_X4 FILLER_10_802 ();
 FILLCELL_X2 FILLER_10_806 ();
 FILLCELL_X1 FILLER_10_808 ();
 FILLCELL_X1 FILLER_10_829 ();
 FILLCELL_X2 FILLER_10_834 ();
 FILLCELL_X2 FILLER_10_856 ();
 FILLCELL_X1 FILLER_10_878 ();
 FILLCELL_X8 FILLER_10_889 ();
 FILLCELL_X2 FILLER_10_897 ();
 FILLCELL_X1 FILLER_10_899 ();
 FILLCELL_X1 FILLER_10_964 ();
 FILLCELL_X1 FILLER_10_972 ();
 FILLCELL_X1 FILLER_10_983 ();
 FILLCELL_X4 FILLER_10_987 ();
 FILLCELL_X2 FILLER_10_991 ();
 FILLCELL_X1 FILLER_10_1016 ();
 FILLCELL_X8 FILLER_10_1021 ();
 FILLCELL_X2 FILLER_10_1029 ();
 FILLCELL_X1 FILLER_10_1031 ();
 FILLCELL_X2 FILLER_10_1044 ();
 FILLCELL_X1 FILLER_10_1046 ();
 FILLCELL_X1 FILLER_10_1081 ();
 FILLCELL_X2 FILLER_10_1103 ();
 FILLCELL_X1 FILLER_10_1113 ();
 FILLCELL_X1 FILLER_10_1121 ();
 FILLCELL_X1 FILLER_10_1126 ();
 FILLCELL_X1 FILLER_10_1131 ();
 FILLCELL_X1 FILLER_10_1136 ();
 FILLCELL_X8 FILLER_10_1140 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_33 ();
 FILLCELL_X4 FILLER_11_41 ();
 FILLCELL_X2 FILLER_11_45 ();
 FILLCELL_X1 FILLER_11_47 ();
 FILLCELL_X1 FILLER_11_68 ();
 FILLCELL_X2 FILLER_11_105 ();
 FILLCELL_X1 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_122 ();
 FILLCELL_X1 FILLER_11_125 ();
 FILLCELL_X2 FILLER_11_134 ();
 FILLCELL_X2 FILLER_11_140 ();
 FILLCELL_X1 FILLER_11_142 ();
 FILLCELL_X8 FILLER_11_187 ();
 FILLCELL_X2 FILLER_11_195 ();
 FILLCELL_X1 FILLER_11_266 ();
 FILLCELL_X1 FILLER_11_307 ();
 FILLCELL_X1 FILLER_11_360 ();
 FILLCELL_X1 FILLER_11_403 ();
 FILLCELL_X2 FILLER_11_455 ();
 FILLCELL_X1 FILLER_11_548 ();
 FILLCELL_X2 FILLER_11_569 ();
 FILLCELL_X1 FILLER_11_571 ();
 FILLCELL_X8 FILLER_11_574 ();
 FILLCELL_X2 FILLER_11_582 ();
 FILLCELL_X1 FILLER_11_630 ();
 FILLCELL_X1 FILLER_11_651 ();
 FILLCELL_X2 FILLER_11_654 ();
 FILLCELL_X1 FILLER_11_656 ();
 FILLCELL_X1 FILLER_11_661 ();
 FILLCELL_X2 FILLER_11_664 ();
 FILLCELL_X4 FILLER_11_676 ();
 FILLCELL_X1 FILLER_11_680 ();
 FILLCELL_X8 FILLER_11_697 ();
 FILLCELL_X4 FILLER_11_705 ();
 FILLCELL_X2 FILLER_11_709 ();
 FILLCELL_X8 FILLER_11_743 ();
 FILLCELL_X4 FILLER_11_751 ();
 FILLCELL_X1 FILLER_11_755 ();
 FILLCELL_X4 FILLER_11_758 ();
 FILLCELL_X4 FILLER_11_764 ();
 FILLCELL_X1 FILLER_11_768 ();
 FILLCELL_X4 FILLER_11_771 ();
 FILLCELL_X2 FILLER_11_775 ();
 FILLCELL_X4 FILLER_11_809 ();
 FILLCELL_X1 FILLER_11_813 ();
 FILLCELL_X4 FILLER_11_816 ();
 FILLCELL_X16 FILLER_11_822 ();
 FILLCELL_X8 FILLER_11_842 ();
 FILLCELL_X2 FILLER_11_850 ();
 FILLCELL_X1 FILLER_11_852 ();
 FILLCELL_X4 FILLER_11_863 ();
 FILLCELL_X1 FILLER_11_867 ();
 FILLCELL_X1 FILLER_11_884 ();
 FILLCELL_X4 FILLER_11_889 ();
 FILLCELL_X1 FILLER_11_893 ();
 FILLCELL_X1 FILLER_11_898 ();
 FILLCELL_X16 FILLER_11_909 ();
 FILLCELL_X4 FILLER_11_925 ();
 FILLCELL_X1 FILLER_11_929 ();
 FILLCELL_X2 FILLER_11_945 ();
 FILLCELL_X1 FILLER_11_947 ();
 FILLCELL_X2 FILLER_11_979 ();
 FILLCELL_X4 FILLER_11_997 ();
 FILLCELL_X1 FILLER_11_1026 ();
 FILLCELL_X4 FILLER_11_1030 ();
 FILLCELL_X2 FILLER_11_1044 ();
 FILLCELL_X1 FILLER_11_1046 ();
 FILLCELL_X2 FILLER_11_1097 ();
 FILLCELL_X2 FILLER_11_1104 ();
 FILLCELL_X2 FILLER_11_1122 ();
 FILLCELL_X1 FILLER_11_1131 ();
 FILLCELL_X4 FILLER_11_1141 ();
 FILLCELL_X2 FILLER_11_1145 ();
 FILLCELL_X1 FILLER_11_1147 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_33 ();
 FILLCELL_X2 FILLER_12_49 ();
 FILLCELL_X1 FILLER_12_51 ();
 FILLCELL_X8 FILLER_12_56 ();
 FILLCELL_X2 FILLER_12_64 ();
 FILLCELL_X1 FILLER_12_66 ();
 FILLCELL_X8 FILLER_12_83 ();
 FILLCELL_X2 FILLER_12_91 ();
 FILLCELL_X1 FILLER_12_95 ();
 FILLCELL_X1 FILLER_12_122 ();
 FILLCELL_X2 FILLER_12_143 ();
 FILLCELL_X2 FILLER_12_149 ();
 FILLCELL_X8 FILLER_12_157 ();
 FILLCELL_X1 FILLER_12_173 ();
 FILLCELL_X1 FILLER_12_194 ();
 FILLCELL_X2 FILLER_12_215 ();
 FILLCELL_X1 FILLER_12_217 ();
 FILLCELL_X4 FILLER_12_278 ();
 FILLCELL_X2 FILLER_12_282 ();
 FILLCELL_X1 FILLER_12_304 ();
 FILLCELL_X1 FILLER_12_360 ();
 FILLCELL_X1 FILLER_12_416 ();
 FILLCELL_X1 FILLER_12_454 ();
 FILLCELL_X2 FILLER_12_535 ();
 FILLCELL_X2 FILLER_12_546 ();
 FILLCELL_X8 FILLER_12_584 ();
 FILLCELL_X4 FILLER_12_595 ();
 FILLCELL_X1 FILLER_12_599 ();
 FILLCELL_X1 FILLER_12_628 ();
 FILLCELL_X1 FILLER_12_632 ();
 FILLCELL_X1 FILLER_12_660 ();
 FILLCELL_X1 FILLER_12_666 ();
 FILLCELL_X8 FILLER_12_669 ();
 FILLCELL_X2 FILLER_12_677 ();
 FILLCELL_X1 FILLER_12_679 ();
 FILLCELL_X1 FILLER_12_684 ();
 FILLCELL_X2 FILLER_12_701 ();
 FILLCELL_X4 FILLER_12_707 ();
 FILLCELL_X2 FILLER_12_711 ();
 FILLCELL_X1 FILLER_12_713 ();
 FILLCELL_X2 FILLER_12_717 ();
 FILLCELL_X2 FILLER_12_723 ();
 FILLCELL_X1 FILLER_12_725 ();
 FILLCELL_X4 FILLER_12_728 ();
 FILLCELL_X2 FILLER_12_735 ();
 FILLCELL_X1 FILLER_12_737 ();
 FILLCELL_X4 FILLER_12_790 ();
 FILLCELL_X1 FILLER_12_794 ();
 FILLCELL_X1 FILLER_12_857 ();
 FILLCELL_X1 FILLER_12_909 ();
 FILLCELL_X2 FILLER_12_1014 ();
 FILLCELL_X4 FILLER_12_1033 ();
 FILLCELL_X2 FILLER_12_1037 ();
 FILLCELL_X1 FILLER_12_1039 ();
 FILLCELL_X1 FILLER_12_1065 ();
 FILLCELL_X1 FILLER_12_1081 ();
 FILLCELL_X1 FILLER_12_1087 ();
 FILLCELL_X2 FILLER_12_1112 ();
 FILLCELL_X2 FILLER_12_1124 ();
 FILLCELL_X8 FILLER_12_1139 ();
 FILLCELL_X1 FILLER_12_1147 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_33 ();
 FILLCELL_X4 FILLER_13_49 ();
 FILLCELL_X2 FILLER_13_87 ();
 FILLCELL_X1 FILLER_13_97 ();
 FILLCELL_X1 FILLER_13_178 ();
 FILLCELL_X1 FILLER_13_181 ();
 FILLCELL_X16 FILLER_13_198 ();
 FILLCELL_X4 FILLER_13_214 ();
 FILLCELL_X2 FILLER_13_218 ();
 FILLCELL_X1 FILLER_13_220 ();
 FILLCELL_X1 FILLER_13_225 ();
 FILLCELL_X1 FILLER_13_230 ();
 FILLCELL_X1 FILLER_13_235 ();
 FILLCELL_X1 FILLER_13_243 ();
 FILLCELL_X4 FILLER_13_250 ();
 FILLCELL_X2 FILLER_13_263 ();
 FILLCELL_X2 FILLER_13_275 ();
 FILLCELL_X1 FILLER_13_287 ();
 FILLCELL_X2 FILLER_13_293 ();
 FILLCELL_X1 FILLER_13_295 ();
 FILLCELL_X2 FILLER_13_305 ();
 FILLCELL_X1 FILLER_13_397 ();
 FILLCELL_X1 FILLER_13_422 ();
 FILLCELL_X1 FILLER_13_446 ();
 FILLCELL_X1 FILLER_13_486 ();
 FILLCELL_X2 FILLER_13_492 ();
 FILLCELL_X1 FILLER_13_494 ();
 FILLCELL_X1 FILLER_13_542 ();
 FILLCELL_X1 FILLER_13_550 ();
 FILLCELL_X2 FILLER_13_578 ();
 FILLCELL_X1 FILLER_13_596 ();
 FILLCELL_X4 FILLER_13_599 ();
 FILLCELL_X2 FILLER_13_603 ();
 FILLCELL_X1 FILLER_13_621 ();
 FILLCELL_X2 FILLER_13_625 ();
 FILLCELL_X4 FILLER_13_671 ();
 FILLCELL_X2 FILLER_13_675 ();
 FILLCELL_X1 FILLER_13_677 ();
 FILLCELL_X4 FILLER_13_686 ();
 FILLCELL_X2 FILLER_13_690 ();
 FILLCELL_X2 FILLER_13_696 ();
 FILLCELL_X4 FILLER_13_752 ();
 FILLCELL_X2 FILLER_13_759 ();
 FILLCELL_X4 FILLER_13_763 ();
 FILLCELL_X2 FILLER_13_783 ();
 FILLCELL_X1 FILLER_13_785 ();
 FILLCELL_X1 FILLER_13_806 ();
 FILLCELL_X2 FILLER_13_809 ();
 FILLCELL_X1 FILLER_13_811 ();
 FILLCELL_X2 FILLER_13_832 ();
 FILLCELL_X2 FILLER_13_853 ();
 FILLCELL_X1 FILLER_13_861 ();
 FILLCELL_X4 FILLER_13_865 ();
 FILLCELL_X2 FILLER_13_869 ();
 FILLCELL_X1 FILLER_13_887 ();
 FILLCELL_X2 FILLER_13_896 ();
 FILLCELL_X1 FILLER_13_898 ();
 FILLCELL_X1 FILLER_13_965 ();
 FILLCELL_X1 FILLER_13_998 ();
 FILLCELL_X1 FILLER_13_1039 ();
 FILLCELL_X1 FILLER_13_1053 ();
 FILLCELL_X2 FILLER_13_1090 ();
 FILLCELL_X8 FILLER_13_1136 ();
 FILLCELL_X4 FILLER_13_1144 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X16 FILLER_14_33 ();
 FILLCELL_X1 FILLER_14_49 ();
 FILLCELL_X4 FILLER_14_66 ();
 FILLCELL_X1 FILLER_14_73 ();
 FILLCELL_X1 FILLER_14_79 ();
 FILLCELL_X4 FILLER_14_104 ();
 FILLCELL_X2 FILLER_14_108 ();
 FILLCELL_X1 FILLER_14_110 ();
 FILLCELL_X1 FILLER_14_115 ();
 FILLCELL_X8 FILLER_14_134 ();
 FILLCELL_X8 FILLER_14_158 ();
 FILLCELL_X2 FILLER_14_166 ();
 FILLCELL_X8 FILLER_14_174 ();
 FILLCELL_X2 FILLER_14_182 ();
 FILLCELL_X2 FILLER_14_186 ();
 FILLCELL_X1 FILLER_14_188 ();
 FILLCELL_X1 FILLER_14_250 ();
 FILLCELL_X1 FILLER_14_265 ();
 FILLCELL_X2 FILLER_14_272 ();
 FILLCELL_X1 FILLER_14_274 ();
 FILLCELL_X2 FILLER_14_293 ();
 FILLCELL_X1 FILLER_14_295 ();
 FILLCELL_X1 FILLER_14_315 ();
 FILLCELL_X2 FILLER_14_323 ();
 FILLCELL_X2 FILLER_14_438 ();
 FILLCELL_X2 FILLER_14_443 ();
 FILLCELL_X2 FILLER_14_486 ();
 FILLCELL_X2 FILLER_14_556 ();
 FILLCELL_X1 FILLER_14_564 ();
 FILLCELL_X1 FILLER_14_585 ();
 FILLCELL_X4 FILLER_14_600 ();
 FILLCELL_X2 FILLER_14_607 ();
 FILLCELL_X4 FILLER_14_611 ();
 FILLCELL_X2 FILLER_14_615 ();
 FILLCELL_X2 FILLER_14_623 ();
 FILLCELL_X1 FILLER_14_625 ();
 FILLCELL_X1 FILLER_14_630 ();
 FILLCELL_X2 FILLER_14_632 ();
 FILLCELL_X1 FILLER_14_656 ();
 FILLCELL_X2 FILLER_14_691 ();
 FILLCELL_X4 FILLER_14_703 ();
 FILLCELL_X2 FILLER_14_707 ();
 FILLCELL_X2 FILLER_14_714 ();
 FILLCELL_X1 FILLER_14_716 ();
 FILLCELL_X1 FILLER_14_736 ();
 FILLCELL_X1 FILLER_14_743 ();
 FILLCELL_X4 FILLER_14_765 ();
 FILLCELL_X1 FILLER_14_769 ();
 FILLCELL_X1 FILLER_14_792 ();
 FILLCELL_X8 FILLER_14_795 ();
 FILLCELL_X1 FILLER_14_803 ();
 FILLCELL_X4 FILLER_14_824 ();
 FILLCELL_X2 FILLER_14_870 ();
 FILLCELL_X1 FILLER_14_879 ();
 FILLCELL_X1 FILLER_14_899 ();
 FILLCELL_X2 FILLER_14_951 ();
 FILLCELL_X2 FILLER_14_973 ();
 FILLCELL_X1 FILLER_14_1062 ();
 FILLCELL_X1 FILLER_14_1067 ();
 FILLCELL_X1 FILLER_14_1097 ();
 FILLCELL_X1 FILLER_14_1111 ();
 FILLCELL_X16 FILLER_14_1132 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X4 FILLER_15_25 ();
 FILLCELL_X16 FILLER_15_36 ();
 FILLCELL_X8 FILLER_15_52 ();
 FILLCELL_X4 FILLER_15_60 ();
 FILLCELL_X2 FILLER_15_64 ();
 FILLCELL_X8 FILLER_15_82 ();
 FILLCELL_X4 FILLER_15_90 ();
 FILLCELL_X1 FILLER_15_94 ();
 FILLCELL_X8 FILLER_15_131 ();
 FILLCELL_X4 FILLER_15_139 ();
 FILLCELL_X2 FILLER_15_143 ();
 FILLCELL_X2 FILLER_15_195 ();
 FILLCELL_X8 FILLER_15_199 ();
 FILLCELL_X2 FILLER_15_207 ();
 FILLCELL_X16 FILLER_15_211 ();
 FILLCELL_X8 FILLER_15_227 ();
 FILLCELL_X1 FILLER_15_265 ();
 FILLCELL_X1 FILLER_15_276 ();
 FILLCELL_X1 FILLER_15_289 ();
 FILLCELL_X1 FILLER_15_296 ();
 FILLCELL_X2 FILLER_15_390 ();
 FILLCELL_X1 FILLER_15_553 ();
 FILLCELL_X1 FILLER_15_571 ();
 FILLCELL_X2 FILLER_15_578 ();
 FILLCELL_X1 FILLER_15_580 ();
 FILLCELL_X8 FILLER_15_583 ();
 FILLCELL_X1 FILLER_15_591 ();
 FILLCELL_X1 FILLER_15_626 ();
 FILLCELL_X2 FILLER_15_637 ();
 FILLCELL_X2 FILLER_15_641 ();
 FILLCELL_X1 FILLER_15_662 ();
 FILLCELL_X8 FILLER_15_677 ();
 FILLCELL_X1 FILLER_15_689 ();
 FILLCELL_X2 FILLER_15_763 ();
 FILLCELL_X1 FILLER_15_765 ();
 FILLCELL_X1 FILLER_15_768 ();
 FILLCELL_X2 FILLER_15_771 ();
 FILLCELL_X2 FILLER_15_813 ();
 FILLCELL_X2 FILLER_15_835 ();
 FILLCELL_X1 FILLER_15_893 ();
 FILLCELL_X2 FILLER_15_926 ();
 FILLCELL_X1 FILLER_15_928 ();
 FILLCELL_X1 FILLER_15_942 ();
 FILLCELL_X2 FILLER_15_1029 ();
 FILLCELL_X1 FILLER_15_1031 ();
 FILLCELL_X4 FILLER_15_1041 ();
 FILLCELL_X1 FILLER_15_1045 ();
 FILLCELL_X1 FILLER_15_1065 ();
 FILLCELL_X16 FILLER_15_1121 ();
 FILLCELL_X8 FILLER_15_1137 ();
 FILLCELL_X2 FILLER_15_1145 ();
 FILLCELL_X1 FILLER_15_1147 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X8 FILLER_16_65 ();
 FILLCELL_X4 FILLER_16_73 ();
 FILLCELL_X2 FILLER_16_77 ();
 FILLCELL_X1 FILLER_16_99 ();
 FILLCELL_X2 FILLER_16_119 ();
 FILLCELL_X1 FILLER_16_121 ();
 FILLCELL_X2 FILLER_16_127 ();
 FILLCELL_X1 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_133 ();
 FILLCELL_X1 FILLER_16_141 ();
 FILLCELL_X2 FILLER_16_160 ();
 FILLCELL_X4 FILLER_16_182 ();
 FILLCELL_X2 FILLER_16_186 ();
 FILLCELL_X4 FILLER_16_204 ();
 FILLCELL_X2 FILLER_16_210 ();
 FILLCELL_X1 FILLER_16_232 ();
 FILLCELL_X1 FILLER_16_243 ();
 FILLCELL_X1 FILLER_16_253 ();
 FILLCELL_X1 FILLER_16_258 ();
 FILLCELL_X1 FILLER_16_286 ();
 FILLCELL_X2 FILLER_16_293 ();
 FILLCELL_X1 FILLER_16_295 ();
 FILLCELL_X1 FILLER_16_299 ();
 FILLCELL_X4 FILLER_16_313 ();
 FILLCELL_X1 FILLER_16_317 ();
 FILLCELL_X1 FILLER_16_353 ();
 FILLCELL_X1 FILLER_16_399 ();
 FILLCELL_X1 FILLER_16_544 ();
 FILLCELL_X2 FILLER_16_566 ();
 FILLCELL_X2 FILLER_16_588 ();
 FILLCELL_X8 FILLER_16_592 ();
 FILLCELL_X1 FILLER_16_600 ();
 FILLCELL_X8 FILLER_16_616 ();
 FILLCELL_X4 FILLER_16_627 ();
 FILLCELL_X1 FILLER_16_635 ();
 FILLCELL_X2 FILLER_16_639 ();
 FILLCELL_X1 FILLER_16_661 ();
 FILLCELL_X2 FILLER_16_664 ();
 FILLCELL_X1 FILLER_16_697 ();
 FILLCELL_X2 FILLER_16_701 ();
 FILLCELL_X4 FILLER_16_707 ();
 FILLCELL_X1 FILLER_16_711 ();
 FILLCELL_X2 FILLER_16_730 ();
 FILLCELL_X4 FILLER_16_734 ();
 FILLCELL_X4 FILLER_16_762 ();
 FILLCELL_X2 FILLER_16_766 ();
 FILLCELL_X1 FILLER_16_768 ();
 FILLCELL_X4 FILLER_16_794 ();
 FILLCELL_X2 FILLER_16_798 ();
 FILLCELL_X2 FILLER_16_829 ();
 FILLCELL_X2 FILLER_16_836 ();
 FILLCELL_X2 FILLER_16_852 ();
 FILLCELL_X1 FILLER_16_854 ();
 FILLCELL_X1 FILLER_16_880 ();
 FILLCELL_X16 FILLER_16_910 ();
 FILLCELL_X1 FILLER_16_936 ();
 FILLCELL_X2 FILLER_16_973 ();
 FILLCELL_X1 FILLER_16_981 ();
 FILLCELL_X1 FILLER_16_985 ();
 FILLCELL_X1 FILLER_16_1029 ();
 FILLCELL_X1 FILLER_16_1041 ();
 FILLCELL_X1 FILLER_16_1068 ();
 FILLCELL_X1 FILLER_16_1072 ();
 FILLCELL_X1 FILLER_16_1076 ();
 FILLCELL_X8 FILLER_16_1135 ();
 FILLCELL_X4 FILLER_16_1143 ();
 FILLCELL_X1 FILLER_16_1147 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_41 ();
 FILLCELL_X1 FILLER_17_45 ();
 FILLCELL_X32 FILLER_17_51 ();
 FILLCELL_X4 FILLER_17_83 ();
 FILLCELL_X1 FILLER_17_87 ();
 FILLCELL_X4 FILLER_17_94 ();
 FILLCELL_X2 FILLER_17_98 ();
 FILLCELL_X1 FILLER_17_146 ();
 FILLCELL_X1 FILLER_17_149 ();
 FILLCELL_X2 FILLER_17_157 ();
 FILLCELL_X2 FILLER_17_167 ();
 FILLCELL_X4 FILLER_17_171 ();
 FILLCELL_X1 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_194 ();
 FILLCELL_X8 FILLER_17_198 ();
 FILLCELL_X4 FILLER_17_206 ();
 FILLCELL_X2 FILLER_17_210 ();
 FILLCELL_X4 FILLER_17_232 ();
 FILLCELL_X2 FILLER_17_236 ();
 FILLCELL_X2 FILLER_17_242 ();
 FILLCELL_X1 FILLER_17_244 ();
 FILLCELL_X1 FILLER_17_248 ();
 FILLCELL_X1 FILLER_17_272 ();
 FILLCELL_X1 FILLER_17_278 ();
 FILLCELL_X1 FILLER_17_281 ();
 FILLCELL_X1 FILLER_17_571 ();
 FILLCELL_X2 FILLER_17_575 ();
 FILLCELL_X2 FILLER_17_597 ();
 FILLCELL_X1 FILLER_17_599 ();
 FILLCELL_X2 FILLER_17_650 ();
 FILLCELL_X2 FILLER_17_684 ();
 FILLCELL_X1 FILLER_17_686 ();
 FILLCELL_X2 FILLER_17_691 ();
 FILLCELL_X1 FILLER_17_693 ();
 FILLCELL_X2 FILLER_17_696 ();
 FILLCELL_X2 FILLER_17_714 ();
 FILLCELL_X1 FILLER_17_716 ();
 FILLCELL_X4 FILLER_17_721 ();
 FILLCELL_X4 FILLER_17_745 ();
 FILLCELL_X2 FILLER_17_749 ();
 FILLCELL_X1 FILLER_17_751 ();
 FILLCELL_X8 FILLER_17_768 ();
 FILLCELL_X4 FILLER_17_776 ();
 FILLCELL_X4 FILLER_17_820 ();
 FILLCELL_X2 FILLER_17_828 ();
 FILLCELL_X1 FILLER_17_834 ();
 FILLCELL_X1 FILLER_17_936 ();
 FILLCELL_X1 FILLER_17_941 ();
 FILLCELL_X1 FILLER_17_953 ();
 FILLCELL_X8 FILLER_17_965 ();
 FILLCELL_X1 FILLER_17_973 ();
 FILLCELL_X1 FILLER_17_997 ();
 FILLCELL_X1 FILLER_17_1008 ();
 FILLCELL_X1 FILLER_17_1012 ();
 FILLCELL_X2 FILLER_17_1049 ();
 FILLCELL_X1 FILLER_17_1055 ();
 FILLCELL_X1 FILLER_17_1115 ();
 FILLCELL_X16 FILLER_17_1129 ();
 FILLCELL_X2 FILLER_17_1145 ();
 FILLCELL_X1 FILLER_17_1147 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X16 FILLER_18_65 ();
 FILLCELL_X1 FILLER_18_81 ();
 FILLCELL_X4 FILLER_18_98 ();
 FILLCELL_X1 FILLER_18_102 ();
 FILLCELL_X2 FILLER_18_127 ();
 FILLCELL_X1 FILLER_18_193 ();
 FILLCELL_X2 FILLER_18_216 ();
 FILLCELL_X1 FILLER_18_218 ();
 FILLCELL_X4 FILLER_18_229 ();
 FILLCELL_X2 FILLER_18_233 ();
 FILLCELL_X2 FILLER_18_245 ();
 FILLCELL_X2 FILLER_18_253 ();
 FILLCELL_X2 FILLER_18_266 ();
 FILLCELL_X1 FILLER_18_273 ();
 FILLCELL_X2 FILLER_18_280 ();
 FILLCELL_X1 FILLER_18_351 ();
 FILLCELL_X2 FILLER_18_454 ();
 FILLCELL_X1 FILLER_18_456 ();
 FILLCELL_X1 FILLER_18_536 ();
 FILLCELL_X4 FILLER_18_549 ();
 FILLCELL_X2 FILLER_18_563 ();
 FILLCELL_X1 FILLER_18_568 ();
 FILLCELL_X4 FILLER_18_576 ();
 FILLCELL_X1 FILLER_18_580 ();
 FILLCELL_X1 FILLER_18_607 ();
 FILLCELL_X8 FILLER_18_610 ();
 FILLCELL_X8 FILLER_18_620 ();
 FILLCELL_X1 FILLER_18_628 ();
 FILLCELL_X4 FILLER_18_664 ();
 FILLCELL_X8 FILLER_18_702 ();
 FILLCELL_X1 FILLER_18_710 ();
 FILLCELL_X16 FILLER_18_715 ();
 FILLCELL_X1 FILLER_18_757 ();
 FILLCELL_X1 FILLER_18_784 ();
 FILLCELL_X4 FILLER_18_865 ();
 FILLCELL_X1 FILLER_18_903 ();
 FILLCELL_X8 FILLER_18_914 ();
 FILLCELL_X2 FILLER_18_922 ();
 FILLCELL_X1 FILLER_18_972 ();
 FILLCELL_X2 FILLER_18_977 ();
 FILLCELL_X1 FILLER_18_979 ();
 FILLCELL_X8 FILLER_18_987 ();
 FILLCELL_X2 FILLER_18_1041 ();
 FILLCELL_X1 FILLER_18_1097 ();
 FILLCELL_X1 FILLER_18_1108 ();
 FILLCELL_X1 FILLER_18_1116 ();
 FILLCELL_X8 FILLER_18_1133 ();
 FILLCELL_X4 FILLER_18_1141 ();
 FILLCELL_X2 FILLER_18_1145 ();
 FILLCELL_X1 FILLER_18_1147 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X8 FILLER_19_17 ();
 FILLCELL_X2 FILLER_19_25 ();
 FILLCELL_X8 FILLER_19_36 ();
 FILLCELL_X2 FILLER_19_44 ();
 FILLCELL_X1 FILLER_19_46 ();
 FILLCELL_X2 FILLER_19_59 ();
 FILLCELL_X2 FILLER_19_91 ();
 FILLCELL_X2 FILLER_19_103 ();
 FILLCELL_X2 FILLER_19_113 ();
 FILLCELL_X1 FILLER_19_115 ();
 FILLCELL_X4 FILLER_19_119 ();
 FILLCELL_X2 FILLER_19_127 ();
 FILLCELL_X1 FILLER_19_129 ();
 FILLCELL_X1 FILLER_19_134 ();
 FILLCELL_X2 FILLER_19_145 ();
 FILLCELL_X1 FILLER_19_147 ();
 FILLCELL_X8 FILLER_19_151 ();
 FILLCELL_X2 FILLER_19_195 ();
 FILLCELL_X1 FILLER_19_197 ();
 FILLCELL_X1 FILLER_19_203 ();
 FILLCELL_X1 FILLER_19_274 ();
 FILLCELL_X4 FILLER_19_300 ();
 FILLCELL_X2 FILLER_19_468 ();
 FILLCELL_X2 FILLER_19_535 ();
 FILLCELL_X1 FILLER_19_537 ();
 FILLCELL_X1 FILLER_19_569 ();
 FILLCELL_X1 FILLER_19_631 ();
 FILLCELL_X8 FILLER_19_650 ();
 FILLCELL_X1 FILLER_19_685 ();
 FILLCELL_X2 FILLER_19_722 ();
 FILLCELL_X8 FILLER_19_752 ();
 FILLCELL_X16 FILLER_19_765 ();
 FILLCELL_X1 FILLER_19_781 ();
 FILLCELL_X2 FILLER_19_802 ();
 FILLCELL_X1 FILLER_19_804 ();
 FILLCELL_X1 FILLER_19_840 ();
 FILLCELL_X4 FILLER_19_921 ();
 FILLCELL_X2 FILLER_19_955 ();
 FILLCELL_X8 FILLER_19_965 ();
 FILLCELL_X1 FILLER_19_973 ();
 FILLCELL_X2 FILLER_19_1027 ();
 FILLCELL_X2 FILLER_19_1065 ();
 FILLCELL_X2 FILLER_19_1123 ();
 FILLCELL_X8 FILLER_19_1133 ();
 FILLCELL_X4 FILLER_19_1141 ();
 FILLCELL_X2 FILLER_19_1145 ();
 FILLCELL_X1 FILLER_19_1147 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_9 ();
 FILLCELL_X2 FILLER_20_13 ();
 FILLCELL_X1 FILLER_20_15 ();
 FILLCELL_X2 FILLER_20_19 ();
 FILLCELL_X1 FILLER_20_21 ();
 FILLCELL_X2 FILLER_20_26 ();
 FILLCELL_X2 FILLER_20_40 ();
 FILLCELL_X1 FILLER_20_60 ();
 FILLCELL_X8 FILLER_20_67 ();
 FILLCELL_X2 FILLER_20_99 ();
 FILLCELL_X1 FILLER_20_101 ();
 FILLCELL_X2 FILLER_20_118 ();
 FILLCELL_X2 FILLER_20_140 ();
 FILLCELL_X1 FILLER_20_158 ();
 FILLCELL_X2 FILLER_20_162 ();
 FILLCELL_X4 FILLER_20_187 ();
 FILLCELL_X1 FILLER_20_225 ();
 FILLCELL_X1 FILLER_20_246 ();
 FILLCELL_X4 FILLER_20_249 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X1 FILLER_20_255 ();
 FILLCELL_X1 FILLER_20_263 ();
 FILLCELL_X1 FILLER_20_467 ();
 FILLCELL_X1 FILLER_20_559 ();
 FILLCELL_X8 FILLER_20_578 ();
 FILLCELL_X1 FILLER_20_586 ();
 FILLCELL_X8 FILLER_20_623 ();
 FILLCELL_X2 FILLER_20_632 ();
 FILLCELL_X1 FILLER_20_634 ();
 FILLCELL_X4 FILLER_20_637 ();
 FILLCELL_X1 FILLER_20_665 ();
 FILLCELL_X2 FILLER_20_686 ();
 FILLCELL_X1 FILLER_20_694 ();
 FILLCELL_X1 FILLER_20_733 ();
 FILLCELL_X16 FILLER_20_738 ();
 FILLCELL_X8 FILLER_20_775 ();
 FILLCELL_X4 FILLER_20_783 ();
 FILLCELL_X8 FILLER_20_807 ();
 FILLCELL_X2 FILLER_20_815 ();
 FILLCELL_X1 FILLER_20_817 ();
 FILLCELL_X2 FILLER_20_821 ();
 FILLCELL_X1 FILLER_20_823 ();
 FILLCELL_X2 FILLER_20_836 ();
 FILLCELL_X2 FILLER_20_878 ();
 FILLCELL_X2 FILLER_20_940 ();
 FILLCELL_X2 FILLER_20_946 ();
 FILLCELL_X2 FILLER_20_970 ();
 FILLCELL_X2 FILLER_20_975 ();
 FILLCELL_X2 FILLER_20_1000 ();
 FILLCELL_X2 FILLER_20_1009 ();
 FILLCELL_X1 FILLER_20_1013 ();
 FILLCELL_X4 FILLER_20_1028 ();
 FILLCELL_X2 FILLER_20_1035 ();
 FILLCELL_X2 FILLER_20_1048 ();
 FILLCELL_X1 FILLER_20_1100 ();
 FILLCELL_X1 FILLER_20_1123 ();
 FILLCELL_X8 FILLER_20_1137 ();
 FILLCELL_X2 FILLER_20_1145 ();
 FILLCELL_X1 FILLER_20_1147 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_15 ();
 FILLCELL_X1 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_30 ();
 FILLCELL_X2 FILLER_21_48 ();
 FILLCELL_X1 FILLER_21_50 ();
 FILLCELL_X2 FILLER_21_53 ();
 FILLCELL_X1 FILLER_21_55 ();
 FILLCELL_X2 FILLER_21_74 ();
 FILLCELL_X1 FILLER_21_76 ();
 FILLCELL_X1 FILLER_21_79 ();
 FILLCELL_X8 FILLER_21_83 ();
 FILLCELL_X1 FILLER_21_91 ();
 FILLCELL_X2 FILLER_21_98 ();
 FILLCELL_X4 FILLER_21_102 ();
 FILLCELL_X2 FILLER_21_106 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X1 FILLER_21_117 ();
 FILLCELL_X4 FILLER_21_120 ();
 FILLCELL_X2 FILLER_21_124 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X2 FILLER_21_140 ();
 FILLCELL_X16 FILLER_21_149 ();
 FILLCELL_X4 FILLER_21_165 ();
 FILLCELL_X1 FILLER_21_169 ();
 FILLCELL_X4 FILLER_21_180 ();
 FILLCELL_X1 FILLER_21_192 ();
 FILLCELL_X1 FILLER_21_209 ();
 FILLCELL_X4 FILLER_21_212 ();
 FILLCELL_X2 FILLER_21_268 ();
 FILLCELL_X1 FILLER_21_282 ();
 FILLCELL_X1 FILLER_21_412 ();
 FILLCELL_X1 FILLER_21_430 ();
 FILLCELL_X1 FILLER_21_436 ();
 FILLCELL_X1 FILLER_21_440 ();
 FILLCELL_X1 FILLER_21_535 ();
 FILLCELL_X2 FILLER_21_540 ();
 FILLCELL_X1 FILLER_21_542 ();
 FILLCELL_X1 FILLER_21_553 ();
 FILLCELL_X1 FILLER_21_575 ();
 FILLCELL_X2 FILLER_21_601 ();
 FILLCELL_X8 FILLER_21_607 ();
 FILLCELL_X4 FILLER_21_615 ();
 FILLCELL_X8 FILLER_21_644 ();
 FILLCELL_X2 FILLER_21_652 ();
 FILLCELL_X1 FILLER_21_660 ();
 FILLCELL_X2 FILLER_21_685 ();
 FILLCELL_X4 FILLER_21_703 ();
 FILLCELL_X2 FILLER_21_710 ();
 FILLCELL_X1 FILLER_21_712 ();
 FILLCELL_X1 FILLER_21_715 ();
 FILLCELL_X4 FILLER_21_719 ();
 FILLCELL_X2 FILLER_21_723 ();
 FILLCELL_X1 FILLER_21_735 ();
 FILLCELL_X1 FILLER_21_756 ();
 FILLCELL_X1 FILLER_21_825 ();
 FILLCELL_X1 FILLER_21_872 ();
 FILLCELL_X8 FILLER_21_883 ();
 FILLCELL_X2 FILLER_21_891 ();
 FILLCELL_X1 FILLER_21_947 ();
 FILLCELL_X2 FILLER_21_962 ();
 FILLCELL_X1 FILLER_21_964 ();
 FILLCELL_X1 FILLER_21_991 ();
 FILLCELL_X1 FILLER_21_996 ();
 FILLCELL_X2 FILLER_21_1025 ();
 FILLCELL_X8 FILLER_21_1046 ();
 FILLCELL_X1 FILLER_21_1054 ();
 FILLCELL_X1 FILLER_21_1064 ();
 FILLCELL_X2 FILLER_21_1068 ();
 FILLCELL_X1 FILLER_21_1070 ();
 FILLCELL_X1 FILLER_21_1073 ();
 FILLCELL_X1 FILLER_21_1130 ();
 FILLCELL_X8 FILLER_21_1133 ();
 FILLCELL_X4 FILLER_21_1141 ();
 FILLCELL_X2 FILLER_21_1145 ();
 FILLCELL_X1 FILLER_21_1147 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_9 ();
 FILLCELL_X1 FILLER_22_35 ();
 FILLCELL_X2 FILLER_22_40 ();
 FILLCELL_X2 FILLER_22_48 ();
 FILLCELL_X4 FILLER_22_56 ();
 FILLCELL_X2 FILLER_22_76 ();
 FILLCELL_X8 FILLER_22_80 ();
 FILLCELL_X1 FILLER_22_100 ();
 FILLCELL_X4 FILLER_22_103 ();
 FILLCELL_X1 FILLER_22_139 ();
 FILLCELL_X2 FILLER_22_156 ();
 FILLCELL_X1 FILLER_22_171 ();
 FILLCELL_X8 FILLER_22_176 ();
 FILLCELL_X1 FILLER_22_184 ();
 FILLCELL_X4 FILLER_22_205 ();
 FILLCELL_X4 FILLER_22_221 ();
 FILLCELL_X2 FILLER_22_265 ();
 FILLCELL_X1 FILLER_22_267 ();
 FILLCELL_X1 FILLER_22_272 ();
 FILLCELL_X2 FILLER_22_293 ();
 FILLCELL_X1 FILLER_22_295 ();
 FILLCELL_X1 FILLER_22_518 ();
 FILLCELL_X2 FILLER_22_537 ();
 FILLCELL_X4 FILLER_22_573 ();
 FILLCELL_X4 FILLER_22_624 ();
 FILLCELL_X2 FILLER_22_628 ();
 FILLCELL_X1 FILLER_22_630 ();
 FILLCELL_X1 FILLER_22_632 ();
 FILLCELL_X8 FILLER_22_676 ();
 FILLCELL_X2 FILLER_22_684 ();
 FILLCELL_X1 FILLER_22_686 ();
 FILLCELL_X8 FILLER_22_689 ();
 FILLCELL_X2 FILLER_22_697 ();
 FILLCELL_X1 FILLER_22_699 ();
 FILLCELL_X4 FILLER_22_702 ();
 FILLCELL_X2 FILLER_22_706 ();
 FILLCELL_X2 FILLER_22_724 ();
 FILLCELL_X1 FILLER_22_726 ();
 FILLCELL_X1 FILLER_22_747 ();
 FILLCELL_X1 FILLER_22_762 ();
 FILLCELL_X8 FILLER_22_773 ();
 FILLCELL_X2 FILLER_22_781 ();
 FILLCELL_X4 FILLER_22_803 ();
 FILLCELL_X1 FILLER_22_844 ();
 FILLCELL_X2 FILLER_22_854 ();
 FILLCELL_X16 FILLER_22_878 ();
 FILLCELL_X2 FILLER_22_894 ();
 FILLCELL_X2 FILLER_22_916 ();
 FILLCELL_X2 FILLER_22_971 ();
 FILLCELL_X2 FILLER_22_1030 ();
 FILLCELL_X1 FILLER_22_1068 ();
 FILLCELL_X2 FILLER_22_1085 ();
 FILLCELL_X1 FILLER_22_1087 ();
 FILLCELL_X8 FILLER_22_1138 ();
 FILLCELL_X2 FILLER_22_1146 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_8 ();
 FILLCELL_X1 FILLER_23_10 ();
 FILLCELL_X4 FILLER_23_63 ();
 FILLCELL_X1 FILLER_23_67 ();
 FILLCELL_X1 FILLER_23_84 ();
 FILLCELL_X4 FILLER_23_119 ();
 FILLCELL_X2 FILLER_23_123 ();
 FILLCELL_X1 FILLER_23_133 ();
 FILLCELL_X1 FILLER_23_136 ();
 FILLCELL_X1 FILLER_23_139 ();
 FILLCELL_X2 FILLER_23_142 ();
 FILLCELL_X1 FILLER_23_148 ();
 FILLCELL_X2 FILLER_23_153 ();
 FILLCELL_X4 FILLER_23_193 ();
 FILLCELL_X2 FILLER_23_197 ();
 FILLCELL_X2 FILLER_23_201 ();
 FILLCELL_X1 FILLER_23_203 ();
 FILLCELL_X4 FILLER_23_252 ();
 FILLCELL_X1 FILLER_23_256 ();
 FILLCELL_X1 FILLER_23_261 ();
 FILLCELL_X1 FILLER_23_266 ();
 FILLCELL_X2 FILLER_23_291 ();
 FILLCELL_X4 FILLER_23_315 ();
 FILLCELL_X2 FILLER_23_399 ();
 FILLCELL_X2 FILLER_23_497 ();
 FILLCELL_X2 FILLER_23_516 ();
 FILLCELL_X1 FILLER_23_540 ();
 FILLCELL_X1 FILLER_23_546 ();
 FILLCELL_X2 FILLER_23_557 ();
 FILLCELL_X1 FILLER_23_566 ();
 FILLCELL_X1 FILLER_23_587 ();
 FILLCELL_X32 FILLER_23_591 ();
 FILLCELL_X8 FILLER_23_623 ();
 FILLCELL_X4 FILLER_23_631 ();
 FILLCELL_X2 FILLER_23_635 ();
 FILLCELL_X1 FILLER_23_637 ();
 FILLCELL_X1 FILLER_23_658 ();
 FILLCELL_X1 FILLER_23_661 ();
 FILLCELL_X1 FILLER_23_675 ();
 FILLCELL_X2 FILLER_23_716 ();
 FILLCELL_X1 FILLER_23_718 ();
 FILLCELL_X4 FILLER_23_775 ();
 FILLCELL_X32 FILLER_23_783 ();
 FILLCELL_X8 FILLER_23_815 ();
 FILLCELL_X4 FILLER_23_823 ();
 FILLCELL_X2 FILLER_23_827 ();
 FILLCELL_X2 FILLER_23_844 ();
 FILLCELL_X1 FILLER_23_846 ();
 FILLCELL_X2 FILLER_23_857 ();
 FILLCELL_X2 FILLER_23_867 ();
 FILLCELL_X1 FILLER_23_869 ();
 FILLCELL_X8 FILLER_23_890 ();
 FILLCELL_X2 FILLER_23_898 ();
 FILLCELL_X1 FILLER_23_970 ();
 FILLCELL_X4 FILLER_23_1007 ();
 FILLCELL_X4 FILLER_23_1043 ();
 FILLCELL_X2 FILLER_23_1047 ();
 FILLCELL_X1 FILLER_23_1088 ();
 FILLCELL_X1 FILLER_23_1100 ();
 FILLCELL_X1 FILLER_23_1130 ();
 FILLCELL_X8 FILLER_23_1136 ();
 FILLCELL_X4 FILLER_23_1144 ();
 FILLCELL_X2 FILLER_24_4 ();
 FILLCELL_X4 FILLER_24_56 ();
 FILLCELL_X2 FILLER_24_60 ();
 FILLCELL_X1 FILLER_24_62 ();
 FILLCELL_X1 FILLER_24_65 ();
 FILLCELL_X1 FILLER_24_73 ();
 FILLCELL_X2 FILLER_24_78 ();
 FILLCELL_X2 FILLER_24_84 ();
 FILLCELL_X2 FILLER_24_102 ();
 FILLCELL_X4 FILLER_24_116 ();
 FILLCELL_X2 FILLER_24_120 ();
 FILLCELL_X4 FILLER_24_124 ();
 FILLCELL_X1 FILLER_24_128 ();
 FILLCELL_X4 FILLER_24_147 ();
 FILLCELL_X1 FILLER_24_189 ();
 FILLCELL_X1 FILLER_24_230 ();
 FILLCELL_X4 FILLER_24_235 ();
 FILLCELL_X1 FILLER_24_239 ();
 FILLCELL_X4 FILLER_24_254 ();
 FILLCELL_X2 FILLER_24_267 ();
 FILLCELL_X1 FILLER_24_269 ();
 FILLCELL_X2 FILLER_24_300 ();
 FILLCELL_X2 FILLER_24_406 ();
 FILLCELL_X2 FILLER_24_542 ();
 FILLCELL_X1 FILLER_24_551 ();
 FILLCELL_X8 FILLER_24_554 ();
 FILLCELL_X4 FILLER_24_562 ();
 FILLCELL_X2 FILLER_24_566 ();
 FILLCELL_X1 FILLER_24_568 ();
 FILLCELL_X4 FILLER_24_598 ();
 FILLCELL_X2 FILLER_24_624 ();
 FILLCELL_X1 FILLER_24_626 ();
 FILLCELL_X2 FILLER_24_682 ();
 FILLCELL_X2 FILLER_24_704 ();
 FILLCELL_X8 FILLER_24_728 ();
 FILLCELL_X4 FILLER_24_736 ();
 FILLCELL_X2 FILLER_24_740 ();
 FILLCELL_X1 FILLER_24_764 ();
 FILLCELL_X1 FILLER_24_767 ();
 FILLCELL_X1 FILLER_24_852 ();
 FILLCELL_X2 FILLER_24_877 ();
 FILLCELL_X1 FILLER_24_898 ();
 FILLCELL_X1 FILLER_24_919 ();
 FILLCELL_X2 FILLER_24_972 ();
 FILLCELL_X8 FILLER_24_1005 ();
 FILLCELL_X4 FILLER_24_1013 ();
 FILLCELL_X2 FILLER_24_1043 ();
 FILLCELL_X4 FILLER_24_1055 ();
 FILLCELL_X1 FILLER_24_1059 ();
 FILLCELL_X1 FILLER_24_1093 ();
 FILLCELL_X16 FILLER_24_1125 ();
 FILLCELL_X4 FILLER_24_1141 ();
 FILLCELL_X2 FILLER_24_1145 ();
 FILLCELL_X1 FILLER_24_1147 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_23 ();
 FILLCELL_X1 FILLER_25_44 ();
 FILLCELL_X1 FILLER_25_64 ();
 FILLCELL_X1 FILLER_25_81 ();
 FILLCELL_X2 FILLER_25_85 ();
 FILLCELL_X4 FILLER_25_91 ();
 FILLCELL_X4 FILLER_25_182 ();
 FILLCELL_X1 FILLER_25_186 ();
 FILLCELL_X4 FILLER_25_203 ();
 FILLCELL_X2 FILLER_25_207 ();
 FILLCELL_X16 FILLER_25_211 ();
 FILLCELL_X2 FILLER_25_227 ();
 FILLCELL_X2 FILLER_25_245 ();
 FILLCELL_X1 FILLER_25_247 ();
 FILLCELL_X1 FILLER_25_253 ();
 FILLCELL_X1 FILLER_25_258 ();
 FILLCELL_X1 FILLER_25_269 ();
 FILLCELL_X1 FILLER_25_310 ();
 FILLCELL_X2 FILLER_25_331 ();
 FILLCELL_X1 FILLER_25_381 ();
 FILLCELL_X1 FILLER_25_394 ();
 FILLCELL_X1 FILLER_25_410 ();
 FILLCELL_X2 FILLER_25_442 ();
 FILLCELL_X1 FILLER_25_489 ();
 FILLCELL_X4 FILLER_25_499 ();
 FILLCELL_X1 FILLER_25_542 ();
 FILLCELL_X1 FILLER_25_550 ();
 FILLCELL_X2 FILLER_25_634 ();
 FILLCELL_X4 FILLER_25_681 ();
 FILLCELL_X2 FILLER_25_691 ();
 FILLCELL_X1 FILLER_25_693 ();
 FILLCELL_X2 FILLER_25_704 ();
 FILLCELL_X1 FILLER_25_753 ();
 FILLCELL_X4 FILLER_25_757 ();
 FILLCELL_X1 FILLER_25_764 ();
 FILLCELL_X4 FILLER_25_770 ();
 FILLCELL_X2 FILLER_25_774 ();
 FILLCELL_X2 FILLER_25_814 ();
 FILLCELL_X2 FILLER_25_825 ();
 FILLCELL_X2 FILLER_25_837 ();
 FILLCELL_X4 FILLER_25_852 ();
 FILLCELL_X1 FILLER_25_856 ();
 FILLCELL_X1 FILLER_25_911 ();
 FILLCELL_X1 FILLER_25_932 ();
 FILLCELL_X1 FILLER_25_942 ();
 FILLCELL_X1 FILLER_25_945 ();
 FILLCELL_X1 FILLER_25_966 ();
 FILLCELL_X1 FILLER_25_971 ();
 FILLCELL_X1 FILLER_25_983 ();
 FILLCELL_X2 FILLER_25_991 ();
 FILLCELL_X2 FILLER_25_1014 ();
 FILLCELL_X1 FILLER_25_1023 ();
 FILLCELL_X2 FILLER_25_1061 ();
 FILLCELL_X1 FILLER_25_1065 ();
 FILLCELL_X1 FILLER_25_1074 ();
 FILLCELL_X1 FILLER_25_1105 ();
 FILLCELL_X16 FILLER_25_1118 ();
 FILLCELL_X8 FILLER_25_1134 ();
 FILLCELL_X4 FILLER_25_1142 ();
 FILLCELL_X2 FILLER_25_1146 ();
 FILLCELL_X4 FILLER_26_1 ();
 FILLCELL_X1 FILLER_26_5 ();
 FILLCELL_X2 FILLER_26_26 ();
 FILLCELL_X1 FILLER_26_28 ();
 FILLCELL_X16 FILLER_26_31 ();
 FILLCELL_X2 FILLER_26_63 ();
 FILLCELL_X1 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_69 ();
 FILLCELL_X2 FILLER_26_73 ();
 FILLCELL_X1 FILLER_26_75 ();
 FILLCELL_X1 FILLER_26_94 ();
 FILLCELL_X1 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_146 ();
 FILLCELL_X2 FILLER_26_158 ();
 FILLCELL_X1 FILLER_26_160 ();
 FILLCELL_X2 FILLER_26_165 ();
 FILLCELL_X1 FILLER_26_167 ();
 FILLCELL_X4 FILLER_26_184 ();
 FILLCELL_X8 FILLER_26_190 ();
 FILLCELL_X4 FILLER_26_198 ();
 FILLCELL_X16 FILLER_26_260 ();
 FILLCELL_X2 FILLER_26_276 ();
 FILLCELL_X1 FILLER_26_278 ();
 FILLCELL_X4 FILLER_26_289 ();
 FILLCELL_X1 FILLER_26_384 ();
 FILLCELL_X1 FILLER_26_430 ();
 FILLCELL_X1 FILLER_26_503 ();
 FILLCELL_X1 FILLER_26_508 ();
 FILLCELL_X1 FILLER_26_519 ();
 FILLCELL_X4 FILLER_26_532 ();
 FILLCELL_X1 FILLER_26_536 ();
 FILLCELL_X1 FILLER_26_557 ();
 FILLCELL_X16 FILLER_26_560 ();
 FILLCELL_X2 FILLER_26_576 ();
 FILLCELL_X2 FILLER_26_584 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X2 FILLER_26_654 ();
 FILLCELL_X1 FILLER_26_656 ();
 FILLCELL_X1 FILLER_26_688 ();
 FILLCELL_X1 FILLER_26_691 ();
 FILLCELL_X1 FILLER_26_710 ();
 FILLCELL_X2 FILLER_26_730 ();
 FILLCELL_X1 FILLER_26_732 ();
 FILLCELL_X2 FILLER_26_755 ();
 FILLCELL_X1 FILLER_26_760 ();
 FILLCELL_X8 FILLER_26_763 ();
 FILLCELL_X2 FILLER_26_799 ();
 FILLCELL_X1 FILLER_26_801 ();
 FILLCELL_X2 FILLER_26_820 ();
 FILLCELL_X1 FILLER_26_838 ();
 FILLCELL_X1 FILLER_26_859 ();
 FILLCELL_X4 FILLER_26_864 ();
 FILLCELL_X2 FILLER_26_868 ();
 FILLCELL_X1 FILLER_26_890 ();
 FILLCELL_X1 FILLER_26_900 ();
 FILLCELL_X1 FILLER_26_903 ();
 FILLCELL_X1 FILLER_26_906 ();
 FILLCELL_X2 FILLER_26_927 ();
 FILLCELL_X2 FILLER_26_1011 ();
 FILLCELL_X1 FILLER_26_1062 ();
 FILLCELL_X1 FILLER_26_1073 ();
 FILLCELL_X1 FILLER_26_1083 ();
 FILLCELL_X4 FILLER_26_1094 ();
 FILLCELL_X2 FILLER_26_1098 ();
 FILLCELL_X1 FILLER_26_1100 ();
 FILLCELL_X2 FILLER_26_1104 ();
 FILLCELL_X1 FILLER_26_1106 ();
 FILLCELL_X16 FILLER_26_1122 ();
 FILLCELL_X8 FILLER_26_1138 ();
 FILLCELL_X2 FILLER_26_1146 ();
 FILLCELL_X4 FILLER_27_45 ();
 FILLCELL_X2 FILLER_27_49 ();
 FILLCELL_X1 FILLER_27_51 ();
 FILLCELL_X4 FILLER_27_86 ();
 FILLCELL_X1 FILLER_27_106 ();
 FILLCELL_X1 FILLER_27_129 ();
 FILLCELL_X8 FILLER_27_133 ();
 FILLCELL_X2 FILLER_27_141 ();
 FILLCELL_X1 FILLER_27_143 ();
 FILLCELL_X4 FILLER_27_164 ();
 FILLCELL_X2 FILLER_27_168 ();
 FILLCELL_X1 FILLER_27_170 ();
 FILLCELL_X8 FILLER_27_173 ();
 FILLCELL_X2 FILLER_27_181 ();
 FILLCELL_X1 FILLER_27_183 ();
 FILLCELL_X8 FILLER_27_231 ();
 FILLCELL_X4 FILLER_27_239 ();
 FILLCELL_X1 FILLER_27_245 ();
 FILLCELL_X1 FILLER_27_389 ();
 FILLCELL_X2 FILLER_27_430 ();
 FILLCELL_X1 FILLER_27_519 ();
 FILLCELL_X1 FILLER_27_525 ();
 FILLCELL_X4 FILLER_27_536 ();
 FILLCELL_X2 FILLER_27_540 ();
 FILLCELL_X2 FILLER_27_592 ();
 FILLCELL_X1 FILLER_27_594 ();
 FILLCELL_X1 FILLER_27_632 ();
 FILLCELL_X4 FILLER_27_648 ();
 FILLCELL_X4 FILLER_27_681 ();
 FILLCELL_X2 FILLER_27_689 ();
 FILLCELL_X2 FILLER_27_724 ();
 FILLCELL_X1 FILLER_27_726 ();
 FILLCELL_X1 FILLER_27_731 ();
 FILLCELL_X2 FILLER_27_752 ();
 FILLCELL_X1 FILLER_27_754 ();
 FILLCELL_X4 FILLER_27_766 ();
 FILLCELL_X1 FILLER_27_784 ();
 FILLCELL_X1 FILLER_27_825 ();
 FILLCELL_X4 FILLER_27_842 ();
 FILLCELL_X2 FILLER_27_846 ();
 FILLCELL_X2 FILLER_27_896 ();
 FILLCELL_X4 FILLER_27_932 ();
 FILLCELL_X2 FILLER_27_936 ();
 FILLCELL_X2 FILLER_27_973 ();
 FILLCELL_X2 FILLER_27_996 ();
 FILLCELL_X4 FILLER_27_1033 ();
 FILLCELL_X1 FILLER_27_1037 ();
 FILLCELL_X4 FILLER_27_1045 ();
 FILLCELL_X2 FILLER_27_1049 ();
 FILLCELL_X8 FILLER_27_1061 ();
 FILLCELL_X2 FILLER_27_1069 ();
 FILLCELL_X32 FILLER_27_1075 ();
 FILLCELL_X32 FILLER_27_1107 ();
 FILLCELL_X8 FILLER_27_1139 ();
 FILLCELL_X1 FILLER_27_1147 ();
 FILLCELL_X8 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_48 ();
 FILLCELL_X1 FILLER_28_72 ();
 FILLCELL_X8 FILLER_28_105 ();
 FILLCELL_X2 FILLER_28_113 ();
 FILLCELL_X1 FILLER_28_115 ();
 FILLCELL_X2 FILLER_28_118 ();
 FILLCELL_X1 FILLER_28_120 ();
 FILLCELL_X4 FILLER_28_214 ();
 FILLCELL_X4 FILLER_28_282 ();
 FILLCELL_X8 FILLER_28_294 ();
 FILLCELL_X2 FILLER_28_302 ();
 FILLCELL_X1 FILLER_28_314 ();
 FILLCELL_X1 FILLER_28_374 ();
 FILLCELL_X1 FILLER_28_379 ();
 FILLCELL_X1 FILLER_28_388 ();
 FILLCELL_X1 FILLER_28_454 ();
 FILLCELL_X8 FILLER_28_541 ();
 FILLCELL_X4 FILLER_28_549 ();
 FILLCELL_X2 FILLER_28_573 ();
 FILLCELL_X2 FILLER_28_581 ();
 FILLCELL_X1 FILLER_28_591 ();
 FILLCELL_X1 FILLER_28_657 ();
 FILLCELL_X1 FILLER_28_683 ();
 FILLCELL_X2 FILLER_28_690 ();
 FILLCELL_X1 FILLER_28_696 ();
 FILLCELL_X2 FILLER_28_720 ();
 FILLCELL_X1 FILLER_28_740 ();
 FILLCELL_X4 FILLER_28_781 ();
 FILLCELL_X1 FILLER_28_787 ();
 FILLCELL_X8 FILLER_28_792 ();
 FILLCELL_X1 FILLER_28_802 ();
 FILLCELL_X1 FILLER_28_805 ();
 FILLCELL_X4 FILLER_28_818 ();
 FILLCELL_X2 FILLER_28_822 ();
 FILLCELL_X4 FILLER_28_844 ();
 FILLCELL_X2 FILLER_28_848 ();
 FILLCELL_X2 FILLER_28_858 ();
 FILLCELL_X1 FILLER_28_860 ();
 FILLCELL_X8 FILLER_28_871 ();
 FILLCELL_X4 FILLER_28_879 ();
 FILLCELL_X1 FILLER_28_883 ();
 FILLCELL_X32 FILLER_28_894 ();
 FILLCELL_X1 FILLER_28_926 ();
 FILLCELL_X1 FILLER_28_947 ();
 FILLCELL_X2 FILLER_28_965 ();
 FILLCELL_X1 FILLER_28_976 ();
 FILLCELL_X1 FILLER_28_982 ();
 FILLCELL_X32 FILLER_28_1011 ();
 FILLCELL_X8 FILLER_28_1043 ();
 FILLCELL_X4 FILLER_28_1051 ();
 FILLCELL_X2 FILLER_28_1055 ();
 FILLCELL_X1 FILLER_28_1057 ();
 FILLCELL_X4 FILLER_28_1065 ();
 FILLCELL_X2 FILLER_28_1069 ();
 FILLCELL_X1 FILLER_28_1071 ();
 FILLCELL_X32 FILLER_28_1087 ();
 FILLCELL_X16 FILLER_28_1119 ();
 FILLCELL_X8 FILLER_28_1135 ();
 FILLCELL_X4 FILLER_28_1143 ();
 FILLCELL_X1 FILLER_28_1147 ();
 FILLCELL_X2 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_3 ();
 FILLCELL_X1 FILLER_29_18 ();
 FILLCELL_X1 FILLER_29_35 ();
 FILLCELL_X1 FILLER_29_38 ();
 FILLCELL_X1 FILLER_29_55 ();
 FILLCELL_X4 FILLER_29_58 ();
 FILLCELL_X2 FILLER_29_64 ();
 FILLCELL_X2 FILLER_29_82 ();
 FILLCELL_X1 FILLER_29_86 ();
 FILLCELL_X2 FILLER_29_97 ();
 FILLCELL_X1 FILLER_29_99 ();
 FILLCELL_X8 FILLER_29_126 ();
 FILLCELL_X2 FILLER_29_154 ();
 FILLCELL_X8 FILLER_29_158 ();
 FILLCELL_X2 FILLER_29_199 ();
 FILLCELL_X1 FILLER_29_206 ();
 FILLCELL_X2 FILLER_29_217 ();
 FILLCELL_X2 FILLER_29_222 ();
 FILLCELL_X1 FILLER_29_224 ();
 FILLCELL_X4 FILLER_29_259 ();
 FILLCELL_X2 FILLER_29_263 ();
 FILLCELL_X1 FILLER_29_265 ();
 FILLCELL_X1 FILLER_29_314 ();
 FILLCELL_X1 FILLER_29_321 ();
 FILLCELL_X2 FILLER_29_328 ();
 FILLCELL_X2 FILLER_29_350 ();
 FILLCELL_X1 FILLER_29_361 ();
 FILLCELL_X1 FILLER_29_369 ();
 FILLCELL_X1 FILLER_29_419 ();
 FILLCELL_X1 FILLER_29_443 ();
 FILLCELL_X1 FILLER_29_447 ();
 FILLCELL_X1 FILLER_29_457 ();
 FILLCELL_X2 FILLER_29_468 ();
 FILLCELL_X1 FILLER_29_470 ();
 FILLCELL_X1 FILLER_29_506 ();
 FILLCELL_X1 FILLER_29_535 ();
 FILLCELL_X2 FILLER_29_601 ();
 FILLCELL_X1 FILLER_29_625 ();
 FILLCELL_X4 FILLER_29_628 ();
 FILLCELL_X2 FILLER_29_672 ();
 FILLCELL_X1 FILLER_29_674 ();
 FILLCELL_X4 FILLER_29_682 ();
 FILLCELL_X1 FILLER_29_696 ();
 FILLCELL_X1 FILLER_29_700 ();
 FILLCELL_X1 FILLER_29_744 ();
 FILLCELL_X1 FILLER_29_749 ();
 FILLCELL_X1 FILLER_29_752 ();
 FILLCELL_X2 FILLER_29_757 ();
 FILLCELL_X8 FILLER_29_775 ();
 FILLCELL_X1 FILLER_29_783 ();
 FILLCELL_X4 FILLER_29_798 ();
 FILLCELL_X1 FILLER_29_828 ();
 FILLCELL_X4 FILLER_29_831 ();
 FILLCELL_X1 FILLER_29_835 ();
 FILLCELL_X4 FILLER_29_860 ();
 FILLCELL_X2 FILLER_29_864 ();
 FILLCELL_X1 FILLER_29_866 ();
 FILLCELL_X1 FILLER_29_885 ();
 FILLCELL_X8 FILLER_29_906 ();
 FILLCELL_X2 FILLER_29_914 ();
 FILLCELL_X1 FILLER_29_916 ();
 FILLCELL_X2 FILLER_29_977 ();
 FILLCELL_X1 FILLER_29_979 ();
 FILLCELL_X16 FILLER_29_982 ();
 FILLCELL_X1 FILLER_29_998 ();
 FILLCELL_X32 FILLER_29_1013 ();
 FILLCELL_X32 FILLER_29_1045 ();
 FILLCELL_X32 FILLER_29_1077 ();
 FILLCELL_X32 FILLER_29_1109 ();
 FILLCELL_X4 FILLER_29_1141 ();
 FILLCELL_X2 FILLER_29_1145 ();
 FILLCELL_X1 FILLER_29_1147 ();
 FILLCELL_X1 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_28 ();
 FILLCELL_X2 FILLER_30_31 ();
 FILLCELL_X1 FILLER_30_33 ();
 FILLCELL_X2 FILLER_30_38 ();
 FILLCELL_X4 FILLER_30_42 ();
 FILLCELL_X2 FILLER_30_46 ();
 FILLCELL_X4 FILLER_30_50 ();
 FILLCELL_X4 FILLER_30_74 ();
 FILLCELL_X2 FILLER_30_78 ();
 FILLCELL_X1 FILLER_30_80 ();
 FILLCELL_X2 FILLER_30_101 ();
 FILLCELL_X2 FILLER_30_107 ();
 FILLCELL_X4 FILLER_30_129 ();
 FILLCELL_X1 FILLER_30_175 ();
 FILLCELL_X1 FILLER_30_181 ();
 FILLCELL_X1 FILLER_30_194 ();
 FILLCELL_X4 FILLER_30_199 ();
 FILLCELL_X2 FILLER_30_203 ();
 FILLCELL_X1 FILLER_30_205 ();
 FILLCELL_X1 FILLER_30_231 ();
 FILLCELL_X4 FILLER_30_247 ();
 FILLCELL_X1 FILLER_30_251 ();
 FILLCELL_X8 FILLER_30_262 ();
 FILLCELL_X2 FILLER_30_270 ();
 FILLCELL_X1 FILLER_30_272 ();
 FILLCELL_X4 FILLER_30_279 ();
 FILLCELL_X1 FILLER_30_283 ();
 FILLCELL_X8 FILLER_30_318 ();
 FILLCELL_X2 FILLER_30_326 ();
 FILLCELL_X1 FILLER_30_350 ();
 FILLCELL_X4 FILLER_30_358 ();
 FILLCELL_X2 FILLER_30_362 ();
 FILLCELL_X2 FILLER_30_371 ();
 FILLCELL_X2 FILLER_30_433 ();
 FILLCELL_X1 FILLER_30_437 ();
 FILLCELL_X1 FILLER_30_505 ();
 FILLCELL_X2 FILLER_30_515 ();
 FILLCELL_X16 FILLER_30_526 ();
 FILLCELL_X4 FILLER_30_542 ();
 FILLCELL_X2 FILLER_30_546 ();
 FILLCELL_X8 FILLER_30_552 ();
 FILLCELL_X1 FILLER_30_562 ();
 FILLCELL_X8 FILLER_30_571 ();
 FILLCELL_X1 FILLER_30_583 ();
 FILLCELL_X2 FILLER_30_600 ();
 FILLCELL_X2 FILLER_30_611 ();
 FILLCELL_X1 FILLER_30_613 ();
 FILLCELL_X2 FILLER_30_618 ();
 FILLCELL_X1 FILLER_30_620 ();
 FILLCELL_X4 FILLER_30_635 ();
 FILLCELL_X1 FILLER_30_650 ();
 FILLCELL_X1 FILLER_30_654 ();
 FILLCELL_X1 FILLER_30_663 ();
 FILLCELL_X8 FILLER_30_668 ();
 FILLCELL_X2 FILLER_30_676 ();
 FILLCELL_X1 FILLER_30_678 ();
 FILLCELL_X1 FILLER_30_685 ();
 FILLCELL_X1 FILLER_30_688 ();
 FILLCELL_X1 FILLER_30_692 ();
 FILLCELL_X1 FILLER_30_696 ();
 FILLCELL_X4 FILLER_30_700 ();
 FILLCELL_X4 FILLER_30_709 ();
 FILLCELL_X1 FILLER_30_713 ();
 FILLCELL_X1 FILLER_30_719 ();
 FILLCELL_X2 FILLER_30_726 ();
 FILLCELL_X2 FILLER_30_731 ();
 FILLCELL_X2 FILLER_30_737 ();
 FILLCELL_X2 FILLER_30_755 ();
 FILLCELL_X1 FILLER_30_757 ();
 FILLCELL_X2 FILLER_30_774 ();
 FILLCELL_X4 FILLER_30_792 ();
 FILLCELL_X2 FILLER_30_796 ();
 FILLCELL_X1 FILLER_30_798 ();
 FILLCELL_X2 FILLER_30_801 ();
 FILLCELL_X1 FILLER_30_803 ();
 FILLCELL_X2 FILLER_30_806 ();
 FILLCELL_X1 FILLER_30_812 ();
 FILLCELL_X1 FILLER_30_831 ();
 FILLCELL_X2 FILLER_30_840 ();
 FILLCELL_X4 FILLER_30_846 ();
 FILLCELL_X2 FILLER_30_882 ();
 FILLCELL_X2 FILLER_30_904 ();
 FILLCELL_X16 FILLER_30_916 ();
 FILLCELL_X8 FILLER_30_932 ();
 FILLCELL_X1 FILLER_30_940 ();
 FILLCELL_X32 FILLER_30_961 ();
 FILLCELL_X32 FILLER_30_993 ();
 FILLCELL_X4 FILLER_30_1025 ();
 FILLCELL_X2 FILLER_30_1029 ();
 FILLCELL_X1 FILLER_30_1031 ();
 FILLCELL_X32 FILLER_30_1052 ();
 FILLCELL_X32 FILLER_30_1084 ();
 FILLCELL_X32 FILLER_30_1116 ();
 FILLCELL_X1 FILLER_31_13 ();
 FILLCELL_X8 FILLER_31_62 ();
 FILLCELL_X1 FILLER_31_70 ();
 FILLCELL_X4 FILLER_31_91 ();
 FILLCELL_X1 FILLER_31_95 ();
 FILLCELL_X2 FILLER_31_164 ();
 FILLCELL_X1 FILLER_31_166 ();
 FILLCELL_X1 FILLER_31_259 ();
 FILLCELL_X1 FILLER_31_264 ();
 FILLCELL_X2 FILLER_31_272 ();
 FILLCELL_X2 FILLER_31_284 ();
 FILLCELL_X1 FILLER_31_302 ();
 FILLCELL_X1 FILLER_31_308 ();
 FILLCELL_X8 FILLER_31_329 ();
 FILLCELL_X4 FILLER_31_337 ();
 FILLCELL_X2 FILLER_31_341 ();
 FILLCELL_X2 FILLER_31_387 ();
 FILLCELL_X1 FILLER_31_398 ();
 FILLCELL_X1 FILLER_31_405 ();
 FILLCELL_X1 FILLER_31_410 ();
 FILLCELL_X1 FILLER_31_428 ();
 FILLCELL_X2 FILLER_31_433 ();
 FILLCELL_X2 FILLER_31_442 ();
 FILLCELL_X1 FILLER_31_451 ();
 FILLCELL_X1 FILLER_31_460 ();
 FILLCELL_X1 FILLER_31_471 ();
 FILLCELL_X1 FILLER_31_476 ();
 FILLCELL_X1 FILLER_31_481 ();
 FILLCELL_X4 FILLER_31_529 ();
 FILLCELL_X2 FILLER_31_533 ();
 FILLCELL_X1 FILLER_31_535 ();
 FILLCELL_X1 FILLER_31_576 ();
 FILLCELL_X2 FILLER_31_581 ();
 FILLCELL_X1 FILLER_31_583 ();
 FILLCELL_X4 FILLER_31_592 ();
 FILLCELL_X4 FILLER_31_600 ();
 FILLCELL_X1 FILLER_31_629 ();
 FILLCELL_X2 FILLER_31_634 ();
 FILLCELL_X1 FILLER_31_636 ();
 FILLCELL_X1 FILLER_31_651 ();
 FILLCELL_X1 FILLER_31_702 ();
 FILLCELL_X4 FILLER_31_716 ();
 FILLCELL_X2 FILLER_31_723 ();
 FILLCELL_X2 FILLER_31_728 ();
 FILLCELL_X1 FILLER_31_730 ();
 FILLCELL_X1 FILLER_31_735 ();
 FILLCELL_X2 FILLER_31_740 ();
 FILLCELL_X1 FILLER_31_742 ();
 FILLCELL_X8 FILLER_31_747 ();
 FILLCELL_X2 FILLER_31_755 ();
 FILLCELL_X1 FILLER_31_757 ();
 FILLCELL_X4 FILLER_31_768 ();
 FILLCELL_X2 FILLER_31_772 ();
 FILLCELL_X1 FILLER_31_792 ();
 FILLCELL_X1 FILLER_31_801 ();
 FILLCELL_X1 FILLER_31_820 ();
 FILLCELL_X1 FILLER_31_853 ();
 FILLCELL_X1 FILLER_31_884 ();
 FILLCELL_X2 FILLER_31_887 ();
 FILLCELL_X1 FILLER_31_889 ();
 FILLCELL_X2 FILLER_31_893 ();
 FILLCELL_X4 FILLER_31_897 ();
 FILLCELL_X1 FILLER_31_901 ();
 FILLCELL_X32 FILLER_31_926 ();
 FILLCELL_X32 FILLER_31_958 ();
 FILLCELL_X32 FILLER_31_990 ();
 FILLCELL_X32 FILLER_31_1022 ();
 FILLCELL_X32 FILLER_31_1054 ();
 FILLCELL_X16 FILLER_31_1086 ();
 FILLCELL_X1 FILLER_31_1102 ();
 FILLCELL_X16 FILLER_31_1123 ();
 FILLCELL_X8 FILLER_31_1139 ();
 FILLCELL_X1 FILLER_31_1147 ();
 FILLCELL_X2 FILLER_32_23 ();
 FILLCELL_X2 FILLER_32_27 ();
 FILLCELL_X2 FILLER_32_32 ();
 FILLCELL_X1 FILLER_32_34 ();
 FILLCELL_X1 FILLER_32_39 ();
 FILLCELL_X1 FILLER_32_44 ();
 FILLCELL_X2 FILLER_32_52 ();
 FILLCELL_X1 FILLER_32_54 ();
 FILLCELL_X1 FILLER_32_71 ();
 FILLCELL_X2 FILLER_32_102 ();
 FILLCELL_X2 FILLER_32_144 ();
 FILLCELL_X1 FILLER_32_157 ();
 FILLCELL_X1 FILLER_32_163 ();
 FILLCELL_X1 FILLER_32_168 ();
 FILLCELL_X1 FILLER_32_175 ();
 FILLCELL_X1 FILLER_32_184 ();
 FILLCELL_X4 FILLER_32_203 ();
 FILLCELL_X1 FILLER_32_211 ();
 FILLCELL_X2 FILLER_32_223 ();
 FILLCELL_X1 FILLER_32_225 ();
 FILLCELL_X2 FILLER_32_263 ();
 FILLCELL_X1 FILLER_32_265 ();
 FILLCELL_X4 FILLER_32_270 ();
 FILLCELL_X1 FILLER_32_274 ();
 FILLCELL_X4 FILLER_32_283 ();
 FILLCELL_X1 FILLER_32_287 ();
 FILLCELL_X1 FILLER_32_308 ();
 FILLCELL_X2 FILLER_32_322 ();
 FILLCELL_X1 FILLER_32_324 ();
 FILLCELL_X1 FILLER_32_347 ();
 FILLCELL_X1 FILLER_32_370 ();
 FILLCELL_X1 FILLER_32_377 ();
 FILLCELL_X8 FILLER_32_412 ();
 FILLCELL_X2 FILLER_32_527 ();
 FILLCELL_X1 FILLER_32_597 ();
 FILLCELL_X2 FILLER_32_614 ();
 FILLCELL_X1 FILLER_32_626 ();
 FILLCELL_X1 FILLER_32_632 ();
 FILLCELL_X4 FILLER_32_647 ();
 FILLCELL_X2 FILLER_32_655 ();
 FILLCELL_X2 FILLER_32_661 ();
 FILLCELL_X1 FILLER_32_663 ();
 FILLCELL_X4 FILLER_32_666 ();
 FILLCELL_X1 FILLER_32_674 ();
 FILLCELL_X1 FILLER_32_679 ();
 FILLCELL_X1 FILLER_32_711 ();
 FILLCELL_X4 FILLER_32_716 ();
 FILLCELL_X2 FILLER_32_724 ();
 FILLCELL_X1 FILLER_32_726 ();
 FILLCELL_X1 FILLER_32_729 ();
 FILLCELL_X2 FILLER_32_746 ();
 FILLCELL_X2 FILLER_32_750 ();
 FILLCELL_X1 FILLER_32_775 ();
 FILLCELL_X1 FILLER_32_778 ();
 FILLCELL_X4 FILLER_32_785 ();
 FILLCELL_X1 FILLER_32_793 ();
 FILLCELL_X2 FILLER_32_798 ();
 FILLCELL_X1 FILLER_32_810 ();
 FILLCELL_X2 FILLER_32_817 ();
 FILLCELL_X1 FILLER_32_819 ();
 FILLCELL_X2 FILLER_32_841 ();
 FILLCELL_X1 FILLER_32_843 ();
 FILLCELL_X2 FILLER_32_860 ();
 FILLCELL_X1 FILLER_32_876 ();
 FILLCELL_X4 FILLER_32_908 ();
 FILLCELL_X1 FILLER_32_912 ();
 FILLCELL_X32 FILLER_32_917 ();
 FILLCELL_X32 FILLER_32_949 ();
 FILLCELL_X8 FILLER_32_981 ();
 FILLCELL_X4 FILLER_32_989 ();
 FILLCELL_X2 FILLER_32_993 ();
 FILLCELL_X32 FILLER_32_1005 ();
 FILLCELL_X32 FILLER_32_1037 ();
 FILLCELL_X32 FILLER_32_1069 ();
 FILLCELL_X16 FILLER_32_1101 ();
 FILLCELL_X4 FILLER_32_1117 ();
 FILLCELL_X1 FILLER_32_1121 ();
 FILLCELL_X16 FILLER_32_1125 ();
 FILLCELL_X4 FILLER_32_1141 ();
 FILLCELL_X2 FILLER_32_1145 ();
 FILLCELL_X1 FILLER_32_1147 ();
 FILLCELL_X1 FILLER_33_21 ();
 FILLCELL_X2 FILLER_33_38 ();
 FILLCELL_X1 FILLER_33_40 ();
 FILLCELL_X2 FILLER_33_61 ();
 FILLCELL_X1 FILLER_33_63 ();
 FILLCELL_X1 FILLER_33_84 ();
 FILLCELL_X8 FILLER_33_96 ();
 FILLCELL_X4 FILLER_33_104 ();
 FILLCELL_X1 FILLER_33_108 ();
 FILLCELL_X8 FILLER_33_113 ();
 FILLCELL_X1 FILLER_33_121 ();
 FILLCELL_X4 FILLER_33_126 ();
 FILLCELL_X4 FILLER_33_134 ();
 FILLCELL_X1 FILLER_33_140 ();
 FILLCELL_X1 FILLER_33_156 ();
 FILLCELL_X1 FILLER_33_164 ();
 FILLCELL_X1 FILLER_33_202 ();
 FILLCELL_X1 FILLER_33_222 ();
 FILLCELL_X1 FILLER_33_227 ();
 FILLCELL_X1 FILLER_33_235 ();
 FILLCELL_X1 FILLER_33_238 ();
 FILLCELL_X2 FILLER_33_242 ();
 FILLCELL_X1 FILLER_33_244 ();
 FILLCELL_X2 FILLER_33_253 ();
 FILLCELL_X1 FILLER_33_255 ();
 FILLCELL_X2 FILLER_33_260 ();
 FILLCELL_X1 FILLER_33_262 ();
 FILLCELL_X4 FILLER_33_285 ();
 FILLCELL_X1 FILLER_33_289 ();
 FILLCELL_X8 FILLER_33_292 ();
 FILLCELL_X8 FILLER_33_360 ();
 FILLCELL_X1 FILLER_33_368 ();
 FILLCELL_X2 FILLER_33_394 ();
 FILLCELL_X1 FILLER_33_396 ();
 FILLCELL_X8 FILLER_33_411 ();
 FILLCELL_X1 FILLER_33_419 ();
 FILLCELL_X2 FILLER_33_430 ();
 FILLCELL_X1 FILLER_33_438 ();
 FILLCELL_X1 FILLER_33_455 ();
 FILLCELL_X2 FILLER_33_491 ();
 FILLCELL_X1 FILLER_33_493 ();
 FILLCELL_X8 FILLER_33_502 ();
 FILLCELL_X2 FILLER_33_510 ();
 FILLCELL_X4 FILLER_33_520 ();
 FILLCELL_X2 FILLER_33_524 ();
 FILLCELL_X1 FILLER_33_526 ();
 FILLCELL_X1 FILLER_33_549 ();
 FILLCELL_X2 FILLER_33_558 ();
 FILLCELL_X1 FILLER_33_560 ();
 FILLCELL_X1 FILLER_33_569 ();
 FILLCELL_X2 FILLER_33_586 ();
 FILLCELL_X2 FILLER_33_604 ();
 FILLCELL_X2 FILLER_33_608 ();
 FILLCELL_X1 FILLER_33_610 ();
 FILLCELL_X2 FILLER_33_631 ();
 FILLCELL_X1 FILLER_33_633 ();
 FILLCELL_X2 FILLER_33_642 ();
 FILLCELL_X1 FILLER_33_664 ();
 FILLCELL_X1 FILLER_33_681 ();
 FILLCELL_X1 FILLER_33_688 ();
 FILLCELL_X8 FILLER_33_692 ();
 FILLCELL_X4 FILLER_33_700 ();
 FILLCELL_X2 FILLER_33_708 ();
 FILLCELL_X1 FILLER_33_710 ();
 FILLCELL_X4 FILLER_33_721 ();
 FILLCELL_X1 FILLER_33_725 ();
 FILLCELL_X2 FILLER_33_730 ();
 FILLCELL_X4 FILLER_33_736 ();
 FILLCELL_X1 FILLER_33_740 ();
 FILLCELL_X2 FILLER_33_755 ();
 FILLCELL_X1 FILLER_33_757 ();
 FILLCELL_X1 FILLER_33_762 ();
 FILLCELL_X2 FILLER_33_767 ();
 FILLCELL_X4 FILLER_33_801 ();
 FILLCELL_X2 FILLER_33_805 ();
 FILLCELL_X8 FILLER_33_834 ();
 FILLCELL_X4 FILLER_33_842 ();
 FILLCELL_X1 FILLER_33_846 ();
 FILLCELL_X4 FILLER_33_881 ();
 FILLCELL_X1 FILLER_33_885 ();
 FILLCELL_X4 FILLER_33_902 ();
 FILLCELL_X32 FILLER_33_928 ();
 FILLCELL_X32 FILLER_33_960 ();
 FILLCELL_X32 FILLER_33_992 ();
 FILLCELL_X32 FILLER_33_1024 ();
 FILLCELL_X32 FILLER_33_1056 ();
 FILLCELL_X32 FILLER_33_1088 ();
 FILLCELL_X16 FILLER_33_1120 ();
 FILLCELL_X8 FILLER_33_1136 ();
 FILLCELL_X4 FILLER_33_1144 ();
 FILLCELL_X2 FILLER_34_1 ();
 FILLCELL_X1 FILLER_34_3 ();
 FILLCELL_X16 FILLER_34_59 ();
 FILLCELL_X2 FILLER_34_75 ();
 FILLCELL_X1 FILLER_34_100 ();
 FILLCELL_X1 FILLER_34_124 ();
 FILLCELL_X2 FILLER_34_189 ();
 FILLCELL_X1 FILLER_34_205 ();
 FILLCELL_X2 FILLER_34_229 ();
 FILLCELL_X8 FILLER_34_242 ();
 FILLCELL_X4 FILLER_34_250 ();
 FILLCELL_X1 FILLER_34_254 ();
 FILLCELL_X1 FILLER_34_258 ();
 FILLCELL_X2 FILLER_34_262 ();
 FILLCELL_X2 FILLER_34_270 ();
 FILLCELL_X4 FILLER_34_300 ();
 FILLCELL_X1 FILLER_34_317 ();
 FILLCELL_X4 FILLER_34_325 ();
 FILLCELL_X1 FILLER_34_329 ();
 FILLCELL_X1 FILLER_34_343 ();
 FILLCELL_X1 FILLER_34_403 ();
 FILLCELL_X1 FILLER_34_431 ();
 FILLCELL_X2 FILLER_34_461 ();
 FILLCELL_X2 FILLER_34_467 ();
 FILLCELL_X1 FILLER_34_472 ();
 FILLCELL_X2 FILLER_34_477 ();
 FILLCELL_X1 FILLER_34_481 ();
 FILLCELL_X1 FILLER_34_484 ();
 FILLCELL_X16 FILLER_34_508 ();
 FILLCELL_X2 FILLER_34_524 ();
 FILLCELL_X2 FILLER_34_546 ();
 FILLCELL_X1 FILLER_34_548 ();
 FILLCELL_X1 FILLER_34_553 ();
 FILLCELL_X4 FILLER_34_558 ();
 FILLCELL_X8 FILLER_34_574 ();
 FILLCELL_X4 FILLER_34_582 ();
 FILLCELL_X1 FILLER_34_588 ();
 FILLCELL_X1 FILLER_34_591 ();
 FILLCELL_X4 FILLER_34_594 ();
 FILLCELL_X1 FILLER_34_602 ();
 FILLCELL_X2 FILLER_34_623 ();
 FILLCELL_X1 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_628 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X1 FILLER_34_651 ();
 FILLCELL_X4 FILLER_34_670 ();
 FILLCELL_X2 FILLER_34_674 ();
 FILLCELL_X1 FILLER_34_676 ();
 FILLCELL_X4 FILLER_34_695 ();
 FILLCELL_X1 FILLER_34_702 ();
 FILLCELL_X1 FILLER_34_719 ();
 FILLCELL_X4 FILLER_34_768 ();
 FILLCELL_X2 FILLER_34_772 ();
 FILLCELL_X1 FILLER_34_774 ();
 FILLCELL_X2 FILLER_34_777 ();
 FILLCELL_X2 FILLER_34_781 ();
 FILLCELL_X1 FILLER_34_783 ();
 FILLCELL_X4 FILLER_34_786 ();
 FILLCELL_X2 FILLER_34_794 ();
 FILLCELL_X1 FILLER_34_796 ();
 FILLCELL_X2 FILLER_34_846 ();
 FILLCELL_X1 FILLER_34_848 ();
 FILLCELL_X8 FILLER_34_851 ();
 FILLCELL_X2 FILLER_34_859 ();
 FILLCELL_X4 FILLER_34_863 ();
 FILLCELL_X4 FILLER_34_869 ();
 FILLCELL_X4 FILLER_34_889 ();
 FILLCELL_X2 FILLER_34_893 ();
 FILLCELL_X1 FILLER_34_895 ();
 FILLCELL_X2 FILLER_34_902 ();
 FILLCELL_X1 FILLER_34_904 ();
 FILLCELL_X32 FILLER_34_925 ();
 FILLCELL_X32 FILLER_34_957 ();
 FILLCELL_X32 FILLER_34_989 ();
 FILLCELL_X32 FILLER_34_1021 ();
 FILLCELL_X32 FILLER_34_1053 ();
 FILLCELL_X32 FILLER_34_1085 ();
 FILLCELL_X16 FILLER_34_1117 ();
 FILLCELL_X8 FILLER_34_1133 ();
 FILLCELL_X4 FILLER_34_1141 ();
 FILLCELL_X2 FILLER_34_1145 ();
 FILLCELL_X1 FILLER_34_1147 ();
 FILLCELL_X4 FILLER_35_37 ();
 FILLCELL_X2 FILLER_35_41 ();
 FILLCELL_X1 FILLER_35_50 ();
 FILLCELL_X2 FILLER_35_53 ();
 FILLCELL_X2 FILLER_35_77 ();
 FILLCELL_X1 FILLER_35_79 ();
 FILLCELL_X2 FILLER_35_119 ();
 FILLCELL_X2 FILLER_35_199 ();
 FILLCELL_X1 FILLER_35_204 ();
 FILLCELL_X4 FILLER_35_211 ();
 FILLCELL_X1 FILLER_35_221 ();
 FILLCELL_X2 FILLER_35_228 ();
 FILLCELL_X4 FILLER_35_233 ();
 FILLCELL_X1 FILLER_35_239 ();
 FILLCELL_X1 FILLER_35_244 ();
 FILLCELL_X1 FILLER_35_250 ();
 FILLCELL_X1 FILLER_35_257 ();
 FILLCELL_X2 FILLER_35_262 ();
 FILLCELL_X1 FILLER_35_264 ();
 FILLCELL_X1 FILLER_35_267 ();
 FILLCELL_X1 FILLER_35_276 ();
 FILLCELL_X1 FILLER_35_286 ();
 FILLCELL_X1 FILLER_35_305 ();
 FILLCELL_X1 FILLER_35_356 ();
 FILLCELL_X2 FILLER_35_380 ();
 FILLCELL_X4 FILLER_35_404 ();
 FILLCELL_X2 FILLER_35_414 ();
 FILLCELL_X1 FILLER_35_443 ();
 FILLCELL_X8 FILLER_35_474 ();
 FILLCELL_X2 FILLER_35_482 ();
 FILLCELL_X1 FILLER_35_484 ();
 FILLCELL_X8 FILLER_35_522 ();
 FILLCELL_X4 FILLER_35_530 ();
 FILLCELL_X1 FILLER_35_534 ();
 FILLCELL_X1 FILLER_35_537 ();
 FILLCELL_X1 FILLER_35_554 ();
 FILLCELL_X1 FILLER_35_559 ();
 FILLCELL_X2 FILLER_35_576 ();
 FILLCELL_X2 FILLER_35_614 ();
 FILLCELL_X1 FILLER_35_616 ();
 FILLCELL_X2 FILLER_35_628 ();
 FILLCELL_X1 FILLER_35_630 ();
 FILLCELL_X1 FILLER_35_635 ();
 FILLCELL_X2 FILLER_35_640 ();
 FILLCELL_X4 FILLER_35_646 ();
 FILLCELL_X2 FILLER_35_650 ();
 FILLCELL_X1 FILLER_35_660 ();
 FILLCELL_X4 FILLER_35_664 ();
 FILLCELL_X1 FILLER_35_668 ();
 FILLCELL_X2 FILLER_35_705 ();
 FILLCELL_X1 FILLER_35_711 ();
 FILLCELL_X1 FILLER_35_716 ();
 FILLCELL_X1 FILLER_35_719 ();
 FILLCELL_X2 FILLER_35_730 ();
 FILLCELL_X4 FILLER_35_736 ();
 FILLCELL_X2 FILLER_35_740 ();
 FILLCELL_X1 FILLER_35_742 ();
 FILLCELL_X1 FILLER_35_759 ();
 FILLCELL_X1 FILLER_35_821 ();
 FILLCELL_X2 FILLER_35_838 ();
 FILLCELL_X1 FILLER_35_840 ();
 FILLCELL_X1 FILLER_35_859 ();
 FILLCELL_X2 FILLER_35_908 ();
 FILLCELL_X1 FILLER_35_910 ();
 FILLCELL_X32 FILLER_35_913 ();
 FILLCELL_X32 FILLER_35_945 ();
 FILLCELL_X32 FILLER_35_977 ();
 FILLCELL_X32 FILLER_35_1009 ();
 FILLCELL_X32 FILLER_35_1041 ();
 FILLCELL_X32 FILLER_35_1073 ();
 FILLCELL_X32 FILLER_35_1105 ();
 FILLCELL_X8 FILLER_35_1137 ();
 FILLCELL_X2 FILLER_35_1145 ();
 FILLCELL_X1 FILLER_35_1147 ();
 FILLCELL_X2 FILLER_36_8 ();
 FILLCELL_X1 FILLER_36_12 ();
 FILLCELL_X1 FILLER_36_15 ();
 FILLCELL_X1 FILLER_36_20 ();
 FILLCELL_X2 FILLER_36_37 ();
 FILLCELL_X4 FILLER_36_44 ();
 FILLCELL_X8 FILLER_36_51 ();
 FILLCELL_X2 FILLER_36_161 ();
 FILLCELL_X16 FILLER_36_167 ();
 FILLCELL_X1 FILLER_36_192 ();
 FILLCELL_X4 FILLER_36_196 ();
 FILLCELL_X2 FILLER_36_213 ();
 FILLCELL_X1 FILLER_36_215 ();
 FILLCELL_X8 FILLER_36_218 ();
 FILLCELL_X2 FILLER_36_226 ();
 FILLCELL_X1 FILLER_36_228 ();
 FILLCELL_X1 FILLER_36_239 ();
 FILLCELL_X1 FILLER_36_245 ();
 FILLCELL_X1 FILLER_36_256 ();
 FILLCELL_X2 FILLER_36_271 ();
 FILLCELL_X1 FILLER_36_273 ();
 FILLCELL_X1 FILLER_36_277 ();
 FILLCELL_X2 FILLER_36_284 ();
 FILLCELL_X2 FILLER_36_297 ();
 FILLCELL_X4 FILLER_36_310 ();
 FILLCELL_X1 FILLER_36_314 ();
 FILLCELL_X8 FILLER_36_322 ();
 FILLCELL_X1 FILLER_36_330 ();
 FILLCELL_X4 FILLER_36_391 ();
 FILLCELL_X2 FILLER_36_442 ();
 FILLCELL_X2 FILLER_36_468 ();
 FILLCELL_X2 FILLER_36_473 ();
 FILLCELL_X1 FILLER_36_482 ();
 FILLCELL_X4 FILLER_36_490 ();
 FILLCELL_X1 FILLER_36_494 ();
 FILLCELL_X1 FILLER_36_505 ();
 FILLCELL_X2 FILLER_36_512 ();
 FILLCELL_X1 FILLER_36_514 ();
 FILLCELL_X16 FILLER_36_531 ();
 FILLCELL_X4 FILLER_36_547 ();
 FILLCELL_X1 FILLER_36_551 ();
 FILLCELL_X8 FILLER_36_596 ();
 FILLCELL_X1 FILLER_36_632 ();
 FILLCELL_X1 FILLER_36_649 ();
 FILLCELL_X4 FILLER_36_666 ();
 FILLCELL_X1 FILLER_36_724 ();
 FILLCELL_X1 FILLER_36_757 ();
 FILLCELL_X2 FILLER_36_781 ();
 FILLCELL_X1 FILLER_36_783 ();
 FILLCELL_X2 FILLER_36_792 ();
 FILLCELL_X1 FILLER_36_794 ();
 FILLCELL_X1 FILLER_36_831 ();
 FILLCELL_X8 FILLER_36_848 ();
 FILLCELL_X4 FILLER_36_856 ();
 FILLCELL_X16 FILLER_36_862 ();
 FILLCELL_X4 FILLER_36_878 ();
 FILLCELL_X2 FILLER_36_882 ();
 FILLCELL_X4 FILLER_36_886 ();
 FILLCELL_X1 FILLER_36_890 ();
 FILLCELL_X32 FILLER_36_931 ();
 FILLCELL_X8 FILLER_36_963 ();
 FILLCELL_X4 FILLER_36_971 ();
 FILLCELL_X2 FILLER_36_975 ();
 FILLCELL_X1 FILLER_36_977 ();
 FILLCELL_X32 FILLER_36_986 ();
 FILLCELL_X1 FILLER_36_1018 ();
 FILLCELL_X1 FILLER_36_1029 ();
 FILLCELL_X32 FILLER_36_1033 ();
 FILLCELL_X32 FILLER_36_1065 ();
 FILLCELL_X1 FILLER_36_1097 ();
 FILLCELL_X16 FILLER_36_1126 ();
 FILLCELL_X2 FILLER_36_1142 ();
 FILLCELL_X1 FILLER_36_1144 ();
 FILLCELL_X4 FILLER_37_70 ();
 FILLCELL_X1 FILLER_37_74 ();
 FILLCELL_X2 FILLER_37_93 ();
 FILLCELL_X4 FILLER_37_115 ();
 FILLCELL_X1 FILLER_37_119 ();
 FILLCELL_X2 FILLER_37_123 ();
 FILLCELL_X1 FILLER_37_141 ();
 FILLCELL_X8 FILLER_37_152 ();
 FILLCELL_X2 FILLER_37_164 ();
 FILLCELL_X1 FILLER_37_170 ();
 FILLCELL_X1 FILLER_37_175 ();
 FILLCELL_X2 FILLER_37_238 ();
 FILLCELL_X4 FILLER_37_246 ();
 FILLCELL_X1 FILLER_37_250 ();
 FILLCELL_X1 FILLER_37_255 ();
 FILLCELL_X1 FILLER_37_278 ();
 FILLCELL_X1 FILLER_37_286 ();
 FILLCELL_X2 FILLER_37_291 ();
 FILLCELL_X1 FILLER_37_293 ();
 FILLCELL_X2 FILLER_37_302 ();
 FILLCELL_X1 FILLER_37_304 ();
 FILLCELL_X1 FILLER_37_312 ();
 FILLCELL_X4 FILLER_37_327 ();
 FILLCELL_X2 FILLER_37_366 ();
 FILLCELL_X1 FILLER_37_368 ();
 FILLCELL_X2 FILLER_37_386 ();
 FILLCELL_X1 FILLER_37_410 ();
 FILLCELL_X1 FILLER_37_433 ();
 FILLCELL_X2 FILLER_37_444 ();
 FILLCELL_X1 FILLER_37_456 ();
 FILLCELL_X1 FILLER_37_461 ();
 FILLCELL_X1 FILLER_37_469 ();
 FILLCELL_X1 FILLER_37_514 ();
 FILLCELL_X1 FILLER_37_521 ();
 FILLCELL_X1 FILLER_37_529 ();
 FILLCELL_X4 FILLER_37_534 ();
 FILLCELL_X2 FILLER_37_538 ();
 FILLCELL_X1 FILLER_37_540 ();
 FILLCELL_X1 FILLER_37_557 ();
 FILLCELL_X2 FILLER_37_574 ();
 FILLCELL_X1 FILLER_37_576 ();
 FILLCELL_X2 FILLER_37_596 ();
 FILLCELL_X4 FILLER_37_635 ();
 FILLCELL_X2 FILLER_37_647 ();
 FILLCELL_X1 FILLER_37_649 ();
 FILLCELL_X2 FILLER_37_662 ();
 FILLCELL_X1 FILLER_37_664 ();
 FILLCELL_X1 FILLER_37_667 ();
 FILLCELL_X8 FILLER_37_671 ();
 FILLCELL_X2 FILLER_37_679 ();
 FILLCELL_X2 FILLER_37_683 ();
 FILLCELL_X8 FILLER_37_693 ();
 FILLCELL_X1 FILLER_37_701 ();
 FILLCELL_X4 FILLER_37_710 ();
 FILLCELL_X2 FILLER_37_714 ();
 FILLCELL_X1 FILLER_37_716 ();
 FILLCELL_X16 FILLER_37_721 ();
 FILLCELL_X4 FILLER_37_737 ();
 FILLCELL_X1 FILLER_37_741 ();
 FILLCELL_X1 FILLER_37_750 ();
 FILLCELL_X8 FILLER_37_754 ();
 FILLCELL_X4 FILLER_37_762 ();
 FILLCELL_X1 FILLER_37_766 ();
 FILLCELL_X2 FILLER_37_780 ();
 FILLCELL_X8 FILLER_37_800 ();
 FILLCELL_X2 FILLER_37_810 ();
 FILLCELL_X1 FILLER_37_812 ();
 FILLCELL_X1 FILLER_37_831 ();
 FILLCELL_X4 FILLER_37_834 ();
 FILLCELL_X1 FILLER_37_838 ();
 FILLCELL_X1 FILLER_37_857 ();
 FILLCELL_X4 FILLER_37_905 ();
 FILLCELL_X1 FILLER_37_914 ();
 FILLCELL_X1 FILLER_37_919 ();
 FILLCELL_X32 FILLER_37_934 ();
 FILLCELL_X8 FILLER_37_966 ();
 FILLCELL_X1 FILLER_37_974 ();
 FILLCELL_X2 FILLER_37_1017 ();
 FILLCELL_X2 FILLER_37_1036 ();
 FILLCELL_X8 FILLER_37_1052 ();
 FILLCELL_X4 FILLER_37_1060 ();
 FILLCELL_X2 FILLER_37_1084 ();
 FILLCELL_X1 FILLER_37_1086 ();
 FILLCELL_X8 FILLER_37_1107 ();
 FILLCELL_X2 FILLER_37_1115 ();
 FILLCELL_X1 FILLER_37_1117 ();
 FILLCELL_X4 FILLER_37_1121 ();
 FILLCELL_X2 FILLER_37_1125 ();
 FILLCELL_X1 FILLER_37_1127 ();
 FILLCELL_X8 FILLER_37_1137 ();
 FILLCELL_X1 FILLER_38_1 ();
 FILLCELL_X8 FILLER_38_46 ();
 FILLCELL_X4 FILLER_38_54 ();
 FILLCELL_X8 FILLER_38_66 ();
 FILLCELL_X2 FILLER_38_74 ();
 FILLCELL_X1 FILLER_38_79 ();
 FILLCELL_X16 FILLER_38_86 ();
 FILLCELL_X4 FILLER_38_109 ();
 FILLCELL_X2 FILLER_38_113 ();
 FILLCELL_X2 FILLER_38_157 ();
 FILLCELL_X2 FILLER_38_185 ();
 FILLCELL_X1 FILLER_38_187 ();
 FILLCELL_X4 FILLER_38_208 ();
 FILLCELL_X1 FILLER_38_244 ();
 FILLCELL_X1 FILLER_38_249 ();
 FILLCELL_X16 FILLER_38_270 ();
 FILLCELL_X2 FILLER_38_286 ();
 FILLCELL_X1 FILLER_38_288 ();
 FILLCELL_X4 FILLER_38_295 ();
 FILLCELL_X1 FILLER_38_299 ();
 FILLCELL_X4 FILLER_38_304 ();
 FILLCELL_X2 FILLER_38_308 ();
 FILLCELL_X4 FILLER_38_316 ();
 FILLCELL_X1 FILLER_38_336 ();
 FILLCELL_X2 FILLER_38_351 ();
 FILLCELL_X2 FILLER_38_357 ();
 FILLCELL_X4 FILLER_38_363 ();
 FILLCELL_X1 FILLER_38_367 ();
 FILLCELL_X2 FILLER_38_420 ();
 FILLCELL_X1 FILLER_38_470 ();
 FILLCELL_X2 FILLER_38_486 ();
 FILLCELL_X1 FILLER_38_488 ();
 FILLCELL_X4 FILLER_38_533 ();
 FILLCELL_X1 FILLER_38_537 ();
 FILLCELL_X4 FILLER_38_564 ();
 FILLCELL_X2 FILLER_38_568 ();
 FILLCELL_X4 FILLER_38_586 ();
 FILLCELL_X1 FILLER_38_590 ();
 FILLCELL_X4 FILLER_38_594 ();
 FILLCELL_X2 FILLER_38_598 ();
 FILLCELL_X1 FILLER_38_600 ();
 FILLCELL_X4 FILLER_38_619 ();
 FILLCELL_X1 FILLER_38_623 ();
 FILLCELL_X2 FILLER_38_626 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X2 FILLER_38_634 ();
 FILLCELL_X1 FILLER_38_640 ();
 FILLCELL_X4 FILLER_38_645 ();
 FILLCELL_X2 FILLER_38_649 ();
 FILLCELL_X1 FILLER_38_667 ();
 FILLCELL_X1 FILLER_38_678 ();
 FILLCELL_X1 FILLER_38_685 ();
 FILLCELL_X2 FILLER_38_718 ();
 FILLCELL_X16 FILLER_38_724 ();
 FILLCELL_X1 FILLER_38_740 ();
 FILLCELL_X2 FILLER_38_757 ();
 FILLCELL_X4 FILLER_38_761 ();
 FILLCELL_X2 FILLER_38_765 ();
 FILLCELL_X1 FILLER_38_787 ();
 FILLCELL_X1 FILLER_38_790 ();
 FILLCELL_X1 FILLER_38_807 ();
 FILLCELL_X1 FILLER_38_824 ();
 FILLCELL_X2 FILLER_38_841 ();
 FILLCELL_X2 FILLER_38_845 ();
 FILLCELL_X1 FILLER_38_867 ();
 FILLCELL_X2 FILLER_38_888 ();
 FILLCELL_X1 FILLER_38_922 ();
 FILLCELL_X32 FILLER_38_925 ();
 FILLCELL_X4 FILLER_38_957 ();
 FILLCELL_X8 FILLER_38_981 ();
 FILLCELL_X4 FILLER_38_989 ();
 FILLCELL_X2 FILLER_38_1013 ();
 FILLCELL_X1 FILLER_38_1026 ();
 FILLCELL_X1 FILLER_38_1040 ();
 FILLCELL_X1 FILLER_38_1069 ();
 FILLCELL_X8 FILLER_38_1080 ();
 FILLCELL_X2 FILLER_38_1088 ();
 FILLCELL_X1 FILLER_38_1090 ();
 FILLCELL_X2 FILLER_38_1137 ();
 FILLCELL_X2 FILLER_39_1 ();
 FILLCELL_X1 FILLER_39_3 ();
 FILLCELL_X2 FILLER_39_9 ();
 FILLCELL_X2 FILLER_39_15 ();
 FILLCELL_X1 FILLER_39_17 ();
 FILLCELL_X2 FILLER_39_51 ();
 FILLCELL_X1 FILLER_39_53 ();
 FILLCELL_X2 FILLER_39_68 ();
 FILLCELL_X2 FILLER_39_88 ();
 FILLCELL_X1 FILLER_39_94 ();
 FILLCELL_X1 FILLER_39_103 ();
 FILLCELL_X2 FILLER_39_119 ();
 FILLCELL_X2 FILLER_39_124 ();
 FILLCELL_X2 FILLER_39_129 ();
 FILLCELL_X2 FILLER_39_134 ();
 FILLCELL_X1 FILLER_39_136 ();
 FILLCELL_X2 FILLER_39_186 ();
 FILLCELL_X1 FILLER_39_188 ();
 FILLCELL_X2 FILLER_39_191 ();
 FILLCELL_X1 FILLER_39_196 ();
 FILLCELL_X16 FILLER_39_199 ();
 FILLCELL_X4 FILLER_39_215 ();
 FILLCELL_X8 FILLER_39_221 ();
 FILLCELL_X2 FILLER_39_237 ();
 FILLCELL_X1 FILLER_39_239 ();
 FILLCELL_X1 FILLER_39_256 ();
 FILLCELL_X16 FILLER_39_293 ();
 FILLCELL_X4 FILLER_39_315 ();
 FILLCELL_X2 FILLER_39_319 ();
 FILLCELL_X1 FILLER_39_326 ();
 FILLCELL_X1 FILLER_39_344 ();
 FILLCELL_X4 FILLER_39_352 ();
 FILLCELL_X1 FILLER_39_387 ();
 FILLCELL_X1 FILLER_39_443 ();
 FILLCELL_X1 FILLER_39_452 ();
 FILLCELL_X1 FILLER_39_458 ();
 FILLCELL_X1 FILLER_39_537 ();
 FILLCELL_X1 FILLER_39_554 ();
 FILLCELL_X2 FILLER_39_557 ();
 FILLCELL_X8 FILLER_39_575 ();
 FILLCELL_X2 FILLER_39_583 ();
 FILLCELL_X1 FILLER_39_585 ();
 FILLCELL_X8 FILLER_39_606 ();
 FILLCELL_X4 FILLER_39_614 ();
 FILLCELL_X1 FILLER_39_668 ();
 FILLCELL_X8 FILLER_39_671 ();
 FILLCELL_X2 FILLER_39_679 ();
 FILLCELL_X8 FILLER_39_699 ();
 FILLCELL_X4 FILLER_39_707 ();
 FILLCELL_X2 FILLER_39_711 ();
 FILLCELL_X1 FILLER_39_731 ();
 FILLCELL_X2 FILLER_39_748 ();
 FILLCELL_X2 FILLER_39_752 ();
 FILLCELL_X4 FILLER_39_770 ();
 FILLCELL_X2 FILLER_39_774 ();
 FILLCELL_X4 FILLER_39_808 ();
 FILLCELL_X1 FILLER_39_812 ();
 FILLCELL_X2 FILLER_39_829 ();
 FILLCELL_X2 FILLER_39_833 ();
 FILLCELL_X16 FILLER_39_855 ();
 FILLCELL_X8 FILLER_39_871 ();
 FILLCELL_X4 FILLER_39_879 ();
 FILLCELL_X1 FILLER_39_898 ();
 FILLCELL_X2 FILLER_39_910 ();
 FILLCELL_X16 FILLER_39_922 ();
 FILLCELL_X8 FILLER_39_938 ();
 FILLCELL_X2 FILLER_39_946 ();
 FILLCELL_X4 FILLER_39_968 ();
 FILLCELL_X2 FILLER_39_1049 ();
 FILLCELL_X1 FILLER_39_1055 ();
 FILLCELL_X16 FILLER_39_1079 ();
 FILLCELL_X1 FILLER_39_1095 ();
 FILLCELL_X2 FILLER_39_1119 ();
 FILLCELL_X1 FILLER_39_1144 ();
 FILLCELL_X1 FILLER_40_1 ();
 FILLCELL_X2 FILLER_40_18 ();
 FILLCELL_X2 FILLER_40_44 ();
 FILLCELL_X2 FILLER_40_48 ();
 FILLCELL_X1 FILLER_40_50 ();
 FILLCELL_X1 FILLER_40_106 ();
 FILLCELL_X1 FILLER_40_111 ();
 FILLCELL_X1 FILLER_40_116 ();
 FILLCELL_X2 FILLER_40_120 ();
 FILLCELL_X1 FILLER_40_122 ();
 FILLCELL_X2 FILLER_40_139 ();
 FILLCELL_X2 FILLER_40_237 ();
 FILLCELL_X1 FILLER_40_239 ();
 FILLCELL_X4 FILLER_40_259 ();
 FILLCELL_X1 FILLER_40_263 ();
 FILLCELL_X4 FILLER_40_268 ();
 FILLCELL_X2 FILLER_40_272 ();
 FILLCELL_X1 FILLER_40_274 ();
 FILLCELL_X4 FILLER_40_315 ();
 FILLCELL_X2 FILLER_40_319 ();
 FILLCELL_X1 FILLER_40_321 ();
 FILLCELL_X1 FILLER_40_340 ();
 FILLCELL_X1 FILLER_40_398 ();
 FILLCELL_X1 FILLER_40_406 ();
 FILLCELL_X1 FILLER_40_414 ();
 FILLCELL_X2 FILLER_40_485 ();
 FILLCELL_X1 FILLER_40_511 ();
 FILLCELL_X2 FILLER_40_538 ();
 FILLCELL_X1 FILLER_40_540 ();
 FILLCELL_X2 FILLER_40_543 ();
 FILLCELL_X2 FILLER_40_612 ();
 FILLCELL_X1 FILLER_40_630 ();
 FILLCELL_X2 FILLER_40_632 ();
 FILLCELL_X1 FILLER_40_696 ();
 FILLCELL_X2 FILLER_40_699 ();
 FILLCELL_X8 FILLER_40_729 ();
 FILLCELL_X2 FILLER_40_737 ();
 FILLCELL_X1 FILLER_40_739 ();
 FILLCELL_X4 FILLER_40_792 ();
 FILLCELL_X1 FILLER_40_796 ();
 FILLCELL_X2 FILLER_40_813 ();
 FILLCELL_X2 FILLER_40_817 ();
 FILLCELL_X1 FILLER_40_819 ();
 FILLCELL_X4 FILLER_40_842 ();
 FILLCELL_X1 FILLER_40_918 ();
 FILLCELL_X32 FILLER_40_922 ();
 FILLCELL_X2 FILLER_40_979 ();
 FILLCELL_X1 FILLER_40_981 ();
 FILLCELL_X2 FILLER_40_1005 ();
 FILLCELL_X1 FILLER_40_1020 ();
 FILLCELL_X2 FILLER_40_1028 ();
 FILLCELL_X1 FILLER_40_1057 ();
 FILLCELL_X1 FILLER_40_1064 ();
 FILLCELL_X1 FILLER_40_1127 ();
 FILLCELL_X2 FILLER_41_4 ();
 FILLCELL_X2 FILLER_41_19 ();
 FILLCELL_X1 FILLER_41_49 ();
 FILLCELL_X4 FILLER_41_55 ();
 FILLCELL_X1 FILLER_41_59 ();
 FILLCELL_X8 FILLER_41_76 ();
 FILLCELL_X2 FILLER_41_84 ();
 FILLCELL_X4 FILLER_41_90 ();
 FILLCELL_X1 FILLER_41_94 ();
 FILLCELL_X1 FILLER_41_116 ();
 FILLCELL_X2 FILLER_41_120 ();
 FILLCELL_X1 FILLER_41_129 ();
 FILLCELL_X4 FILLER_41_134 ();
 FILLCELL_X2 FILLER_41_138 ();
 FILLCELL_X1 FILLER_41_144 ();
 FILLCELL_X4 FILLER_41_153 ();
 FILLCELL_X1 FILLER_41_157 ();
 FILLCELL_X2 FILLER_41_165 ();
 FILLCELL_X4 FILLER_41_175 ();
 FILLCELL_X2 FILLER_41_179 ();
 FILLCELL_X4 FILLER_41_200 ();
 FILLCELL_X2 FILLER_41_204 ();
 FILLCELL_X8 FILLER_41_218 ();
 FILLCELL_X4 FILLER_41_232 ();
 FILLCELL_X2 FILLER_41_236 ();
 FILLCELL_X1 FILLER_41_238 ();
 FILLCELL_X1 FILLER_41_247 ();
 FILLCELL_X1 FILLER_41_270 ();
 FILLCELL_X4 FILLER_41_273 ();
 FILLCELL_X2 FILLER_41_277 ();
 FILLCELL_X1 FILLER_41_279 ();
 FILLCELL_X2 FILLER_41_300 ();
 FILLCELL_X1 FILLER_41_302 ();
 FILLCELL_X4 FILLER_41_305 ();
 FILLCELL_X1 FILLER_41_309 ();
 FILLCELL_X1 FILLER_41_330 ();
 FILLCELL_X1 FILLER_41_333 ();
 FILLCELL_X1 FILLER_41_356 ();
 FILLCELL_X2 FILLER_41_371 ();
 FILLCELL_X2 FILLER_41_375 ();
 FILLCELL_X2 FILLER_41_428 ();
 FILLCELL_X1 FILLER_41_474 ();
 FILLCELL_X2 FILLER_41_480 ();
 FILLCELL_X2 FILLER_41_489 ();
 FILLCELL_X1 FILLER_41_533 ();
 FILLCELL_X2 FILLER_41_550 ();
 FILLCELL_X1 FILLER_41_552 ();
 FILLCELL_X2 FILLER_41_577 ();
 FILLCELL_X4 FILLER_41_601 ();
 FILLCELL_X2 FILLER_41_605 ();
 FILLCELL_X1 FILLER_41_607 ();
 FILLCELL_X4 FILLER_41_613 ();
 FILLCELL_X2 FILLER_41_617 ();
 FILLCELL_X2 FILLER_41_635 ();
 FILLCELL_X1 FILLER_41_655 ();
 FILLCELL_X1 FILLER_41_658 ();
 FILLCELL_X4 FILLER_41_677 ();
 FILLCELL_X2 FILLER_41_681 ();
 FILLCELL_X1 FILLER_41_683 ();
 FILLCELL_X1 FILLER_41_686 ();
 FILLCELL_X4 FILLER_41_719 ();
 FILLCELL_X1 FILLER_41_723 ();
 FILLCELL_X1 FILLER_41_732 ();
 FILLCELL_X1 FILLER_41_749 ();
 FILLCELL_X1 FILLER_41_753 ();
 FILLCELL_X1 FILLER_41_757 ();
 FILLCELL_X1 FILLER_41_761 ();
 FILLCELL_X1 FILLER_41_765 ();
 FILLCELL_X1 FILLER_41_782 ();
 FILLCELL_X2 FILLER_41_801 ();
 FILLCELL_X1 FILLER_41_803 ();
 FILLCELL_X2 FILLER_41_824 ();
 FILLCELL_X8 FILLER_41_828 ();
 FILLCELL_X2 FILLER_41_903 ();
 FILLCELL_X1 FILLER_41_905 ();
 FILLCELL_X8 FILLER_41_919 ();
 FILLCELL_X2 FILLER_41_927 ();
 FILLCELL_X4 FILLER_41_949 ();
 FILLCELL_X2 FILLER_41_953 ();
 FILLCELL_X1 FILLER_41_955 ();
 FILLCELL_X2 FILLER_41_986 ();
 FILLCELL_X1 FILLER_41_995 ();
 FILLCELL_X1 FILLER_41_1018 ();
 FILLCELL_X2 FILLER_41_1037 ();
 FILLCELL_X1 FILLER_41_1053 ();
 FILLCELL_X2 FILLER_41_1064 ();
 FILLCELL_X16 FILLER_41_1082 ();
 FILLCELL_X1 FILLER_41_1111 ();
 FILLCELL_X1 FILLER_41_1115 ();
 FILLCELL_X2 FILLER_42_1 ();
 FILLCELL_X1 FILLER_42_3 ();
 FILLCELL_X2 FILLER_42_24 ();
 FILLCELL_X4 FILLER_42_62 ();
 FILLCELL_X2 FILLER_42_66 ();
 FILLCELL_X2 FILLER_42_76 ();
 FILLCELL_X1 FILLER_42_112 ();
 FILLCELL_X8 FILLER_42_129 ();
 FILLCELL_X2 FILLER_42_137 ();
 FILLCELL_X2 FILLER_42_141 ();
 FILLCELL_X2 FILLER_42_190 ();
 FILLCELL_X1 FILLER_42_192 ();
 FILLCELL_X4 FILLER_42_195 ();
 FILLCELL_X1 FILLER_42_199 ();
 FILLCELL_X2 FILLER_42_202 ();
 FILLCELL_X2 FILLER_42_242 ();
 FILLCELL_X2 FILLER_42_254 ();
 FILLCELL_X1 FILLER_42_256 ();
 FILLCELL_X1 FILLER_42_297 ();
 FILLCELL_X8 FILLER_42_318 ();
 FILLCELL_X1 FILLER_42_340 ();
 FILLCELL_X2 FILLER_42_346 ();
 FILLCELL_X2 FILLER_42_377 ();
 FILLCELL_X1 FILLER_42_379 ();
 FILLCELL_X2 FILLER_42_429 ();
 FILLCELL_X1 FILLER_42_476 ();
 FILLCELL_X1 FILLER_42_531 ();
 FILLCELL_X16 FILLER_42_552 ();
 FILLCELL_X4 FILLER_42_568 ();
 FILLCELL_X4 FILLER_42_590 ();
 FILLCELL_X2 FILLER_42_594 ();
 FILLCELL_X1 FILLER_42_596 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X8 FILLER_42_632 ();
 FILLCELL_X1 FILLER_42_640 ();
 FILLCELL_X4 FILLER_42_697 ();
 FILLCELL_X2 FILLER_42_701 ();
 FILLCELL_X1 FILLER_42_703 ();
 FILLCELL_X1 FILLER_42_720 ();
 FILLCELL_X1 FILLER_42_749 ();
 FILLCELL_X8 FILLER_42_768 ();
 FILLCELL_X4 FILLER_42_776 ();
 FILLCELL_X2 FILLER_42_780 ();
 FILLCELL_X8 FILLER_42_815 ();
 FILLCELL_X1 FILLER_42_823 ();
 FILLCELL_X2 FILLER_42_869 ();
 FILLCELL_X1 FILLER_42_871 ();
 FILLCELL_X2 FILLER_42_877 ();
 FILLCELL_X1 FILLER_42_895 ();
 FILLCELL_X2 FILLER_42_913 ();
 FILLCELL_X4 FILLER_42_935 ();
 FILLCELL_X2 FILLER_42_939 ();
 FILLCELL_X1 FILLER_42_964 ();
 FILLCELL_X1 FILLER_42_975 ();
 FILLCELL_X1 FILLER_42_990 ();
 FILLCELL_X1 FILLER_42_995 ();
 FILLCELL_X1 FILLER_42_1001 ();
 FILLCELL_X2 FILLER_42_1047 ();
 FILLCELL_X1 FILLER_42_1060 ();
 FILLCELL_X8 FILLER_42_1075 ();
 FILLCELL_X1 FILLER_42_1098 ();
 FILLCELL_X1 FILLER_42_1127 ();
 FILLCELL_X4 FILLER_43_1 ();
 FILLCELL_X2 FILLER_43_5 ();
 FILLCELL_X2 FILLER_43_39 ();
 FILLCELL_X4 FILLER_43_57 ();
 FILLCELL_X8 FILLER_43_79 ();
 FILLCELL_X2 FILLER_43_87 ();
 FILLCELL_X1 FILLER_43_89 ();
 FILLCELL_X2 FILLER_43_92 ();
 FILLCELL_X1 FILLER_43_94 ();
 FILLCELL_X1 FILLER_43_97 ();
 FILLCELL_X4 FILLER_43_117 ();
 FILLCELL_X2 FILLER_43_124 ();
 FILLCELL_X1 FILLER_43_126 ();
 FILLCELL_X1 FILLER_43_131 ();
 FILLCELL_X8 FILLER_43_156 ();
 FILLCELL_X1 FILLER_43_164 ();
 FILLCELL_X4 FILLER_43_169 ();
 FILLCELL_X1 FILLER_43_173 ();
 FILLCELL_X2 FILLER_43_206 ();
 FILLCELL_X2 FILLER_43_226 ();
 FILLCELL_X1 FILLER_43_228 ();
 FILLCELL_X2 FILLER_43_311 ();
 FILLCELL_X8 FILLER_43_323 ();
 FILLCELL_X1 FILLER_43_331 ();
 FILLCELL_X1 FILLER_43_362 ();
 FILLCELL_X4 FILLER_43_387 ();
 FILLCELL_X2 FILLER_43_404 ();
 FILLCELL_X1 FILLER_43_406 ();
 FILLCELL_X1 FILLER_43_568 ();
 FILLCELL_X1 FILLER_43_571 ();
 FILLCELL_X1 FILLER_43_574 ();
 FILLCELL_X1 FILLER_43_579 ();
 FILLCELL_X16 FILLER_43_614 ();
 FILLCELL_X2 FILLER_43_646 ();
 FILLCELL_X4 FILLER_43_650 ();
 FILLCELL_X2 FILLER_43_654 ();
 FILLCELL_X8 FILLER_43_658 ();
 FILLCELL_X2 FILLER_43_688 ();
 FILLCELL_X1 FILLER_43_690 ();
 FILLCELL_X1 FILLER_43_701 ();
 FILLCELL_X2 FILLER_43_722 ();
 FILLCELL_X1 FILLER_43_724 ();
 FILLCELL_X1 FILLER_43_747 ();
 FILLCELL_X1 FILLER_43_826 ();
 FILLCELL_X2 FILLER_43_837 ();
 FILLCELL_X1 FILLER_43_847 ();
 FILLCELL_X4 FILLER_43_879 ();
 FILLCELL_X1 FILLER_43_883 ();
 FILLCELL_X4 FILLER_43_899 ();
 FILLCELL_X1 FILLER_43_903 ();
 FILLCELL_X8 FILLER_43_915 ();
 FILLCELL_X4 FILLER_43_923 ();
 FILLCELL_X2 FILLER_43_927 ();
 FILLCELL_X1 FILLER_43_929 ();
 FILLCELL_X16 FILLER_43_937 ();
 FILLCELL_X2 FILLER_43_953 ();
 FILLCELL_X8 FILLER_43_970 ();
 FILLCELL_X2 FILLER_43_978 ();
 FILLCELL_X1 FILLER_43_980 ();
 FILLCELL_X2 FILLER_43_986 ();
 FILLCELL_X1 FILLER_43_988 ();
 FILLCELL_X2 FILLER_43_1049 ();
 FILLCELL_X1 FILLER_43_1064 ();
 FILLCELL_X2 FILLER_43_1083 ();
 FILLCELL_X2 FILLER_43_1109 ();
 FILLCELL_X2 FILLER_44_11 ();
 FILLCELL_X2 FILLER_44_33 ();
 FILLCELL_X4 FILLER_44_223 ();
 FILLCELL_X1 FILLER_44_259 ();
 FILLCELL_X2 FILLER_44_264 ();
 FILLCELL_X1 FILLER_44_270 ();
 FILLCELL_X1 FILLER_44_275 ();
 FILLCELL_X1 FILLER_44_306 ();
 FILLCELL_X2 FILLER_44_320 ();
 FILLCELL_X1 FILLER_44_360 ();
 FILLCELL_X1 FILLER_44_385 ();
 FILLCELL_X1 FILLER_44_410 ();
 FILLCELL_X4 FILLER_44_475 ();
 FILLCELL_X1 FILLER_44_501 ();
 FILLCELL_X1 FILLER_44_525 ();
 FILLCELL_X1 FILLER_44_547 ();
 FILLCELL_X2 FILLER_44_605 ();
 FILLCELL_X1 FILLER_44_632 ();
 FILLCELL_X8 FILLER_44_635 ();
 FILLCELL_X2 FILLER_44_643 ();
 FILLCELL_X2 FILLER_44_647 ();
 FILLCELL_X2 FILLER_44_676 ();
 FILLCELL_X8 FILLER_44_703 ();
 FILLCELL_X4 FILLER_44_711 ();
 FILLCELL_X2 FILLER_44_715 ();
 FILLCELL_X1 FILLER_44_717 ();
 FILLCELL_X8 FILLER_44_738 ();
 FILLCELL_X4 FILLER_44_746 ();
 FILLCELL_X2 FILLER_44_750 ();
 FILLCELL_X1 FILLER_44_752 ();
 FILLCELL_X4 FILLER_44_818 ();
 FILLCELL_X2 FILLER_44_822 ();
 FILLCELL_X1 FILLER_44_824 ();
 FILLCELL_X4 FILLER_44_835 ();
 FILLCELL_X2 FILLER_44_869 ();
 FILLCELL_X1 FILLER_44_881 ();
 FILLCELL_X1 FILLER_44_893 ();
 FILLCELL_X1 FILLER_44_903 ();
 FILLCELL_X8 FILLER_44_911 ();
 FILLCELL_X4 FILLER_44_919 ();
 FILLCELL_X4 FILLER_44_979 ();
 FILLCELL_X2 FILLER_44_1026 ();
 FILLCELL_X2 FILLER_44_1054 ();
 FILLCELL_X1 FILLER_44_1056 ();
 FILLCELL_X1 FILLER_44_1083 ();
 FILLCELL_X1 FILLER_44_1088 ();
 FILLCELL_X1 FILLER_44_1103 ();
 FILLCELL_X2 FILLER_44_1110 ();
 FILLCELL_X2 FILLER_44_1146 ();
 FILLCELL_X1 FILLER_45_3 ();
 FILLCELL_X1 FILLER_45_20 ();
 FILLCELL_X1 FILLER_45_53 ();
 FILLCELL_X4 FILLER_45_86 ();
 FILLCELL_X2 FILLER_45_90 ();
 FILLCELL_X1 FILLER_45_92 ();
 FILLCELL_X4 FILLER_45_96 ();
 FILLCELL_X2 FILLER_45_100 ();
 FILLCELL_X1 FILLER_45_102 ();
 FILLCELL_X8 FILLER_45_110 ();
 FILLCELL_X4 FILLER_45_118 ();
 FILLCELL_X2 FILLER_45_122 ();
 FILLCELL_X1 FILLER_45_152 ();
 FILLCELL_X2 FILLER_45_169 ();
 FILLCELL_X1 FILLER_45_187 ();
 FILLCELL_X2 FILLER_45_204 ();
 FILLCELL_X1 FILLER_45_222 ();
 FILLCELL_X1 FILLER_45_227 ();
 FILLCELL_X4 FILLER_45_238 ();
 FILLCELL_X1 FILLER_45_245 ();
 FILLCELL_X2 FILLER_45_264 ();
 FILLCELL_X1 FILLER_45_266 ();
 FILLCELL_X2 FILLER_45_294 ();
 FILLCELL_X2 FILLER_45_312 ();
 FILLCELL_X1 FILLER_45_314 ();
 FILLCELL_X4 FILLER_45_318 ();
 FILLCELL_X2 FILLER_45_322 ();
 FILLCELL_X1 FILLER_45_324 ();
 FILLCELL_X1 FILLER_45_366 ();
 FILLCELL_X2 FILLER_45_490 ();
 FILLCELL_X4 FILLER_45_624 ();
 FILLCELL_X16 FILLER_45_728 ();
 FILLCELL_X2 FILLER_45_744 ();
 FILLCELL_X2 FILLER_45_821 ();
 FILLCELL_X4 FILLER_45_827 ();
 FILLCELL_X2 FILLER_45_831 ();
 FILLCELL_X1 FILLER_45_833 ();
 FILLCELL_X4 FILLER_45_838 ();
 FILLCELL_X2 FILLER_45_842 ();
 FILLCELL_X2 FILLER_45_847 ();
 FILLCELL_X1 FILLER_45_849 ();
 FILLCELL_X4 FILLER_45_891 ();
 FILLCELL_X16 FILLER_45_918 ();
 FILLCELL_X2 FILLER_45_951 ();
 FILLCELL_X1 FILLER_45_953 ();
 FILLCELL_X1 FILLER_45_960 ();
 FILLCELL_X1 FILLER_45_968 ();
 FILLCELL_X2 FILLER_45_979 ();
 FILLCELL_X2 FILLER_45_1024 ();
 FILLCELL_X1 FILLER_45_1029 ();
 FILLCELL_X1 FILLER_45_1034 ();
 FILLCELL_X1 FILLER_45_1039 ();
 FILLCELL_X1 FILLER_45_1047 ();
 FILLCELL_X1 FILLER_45_1057 ();
 FILLCELL_X2 FILLER_45_1071 ();
 FILLCELL_X2 FILLER_45_1110 ();
 FILLCELL_X1 FILLER_45_1112 ();
 FILLCELL_X1 FILLER_45_1127 ();
 FILLCELL_X1 FILLER_45_1131 ();
 FILLCELL_X1 FILLER_45_1142 ();
 FILLCELL_X2 FILLER_46_4 ();
 FILLCELL_X1 FILLER_46_10 ();
 FILLCELL_X1 FILLER_46_47 ();
 FILLCELL_X16 FILLER_46_64 ();
 FILLCELL_X4 FILLER_46_80 ();
 FILLCELL_X1 FILLER_46_84 ();
 FILLCELL_X1 FILLER_46_101 ();
 FILLCELL_X1 FILLER_46_106 ();
 FILLCELL_X1 FILLER_46_115 ();
 FILLCELL_X2 FILLER_46_132 ();
 FILLCELL_X2 FILLER_46_156 ();
 FILLCELL_X1 FILLER_46_158 ();
 FILLCELL_X16 FILLER_46_180 ();
 FILLCELL_X8 FILLER_46_198 ();
 FILLCELL_X16 FILLER_46_214 ();
 FILLCELL_X1 FILLER_46_230 ();
 FILLCELL_X2 FILLER_46_235 ();
 FILLCELL_X4 FILLER_46_241 ();
 FILLCELL_X2 FILLER_46_245 ();
 FILLCELL_X8 FILLER_46_250 ();
 FILLCELL_X1 FILLER_46_258 ();
 FILLCELL_X1 FILLER_46_263 ();
 FILLCELL_X1 FILLER_46_284 ();
 FILLCELL_X1 FILLER_46_305 ();
 FILLCELL_X4 FILLER_46_334 ();
 FILLCELL_X1 FILLER_46_368 ();
 FILLCELL_X2 FILLER_46_383 ();
 FILLCELL_X2 FILLER_46_420 ();
 FILLCELL_X1 FILLER_46_422 ();
 FILLCELL_X4 FILLER_46_548 ();
 FILLCELL_X1 FILLER_46_552 ();
 FILLCELL_X2 FILLER_46_571 ();
 FILLCELL_X1 FILLER_46_609 ();
 FILLCELL_X1 FILLER_46_630 ();
 FILLCELL_X8 FILLER_46_634 ();
 FILLCELL_X2 FILLER_46_642 ();
 FILLCELL_X1 FILLER_46_644 ();
 FILLCELL_X4 FILLER_46_665 ();
 FILLCELL_X2 FILLER_46_669 ();
 FILLCELL_X1 FILLER_46_671 ();
 FILLCELL_X2 FILLER_46_682 ();
 FILLCELL_X1 FILLER_46_694 ();
 FILLCELL_X1 FILLER_46_699 ();
 FILLCELL_X2 FILLER_46_712 ();
 FILLCELL_X2 FILLER_46_724 ();
 FILLCELL_X1 FILLER_46_726 ();
 FILLCELL_X2 FILLER_46_747 ();
 FILLCELL_X1 FILLER_46_749 ();
 FILLCELL_X8 FILLER_46_752 ();
 FILLCELL_X4 FILLER_46_794 ();
 FILLCELL_X8 FILLER_46_818 ();
 FILLCELL_X1 FILLER_46_826 ();
 FILLCELL_X2 FILLER_46_875 ();
 FILLCELL_X1 FILLER_46_895 ();
 FILLCELL_X1 FILLER_46_902 ();
 FILLCELL_X1 FILLER_46_913 ();
 FILLCELL_X2 FILLER_46_916 ();
 FILLCELL_X1 FILLER_46_975 ();
 FILLCELL_X4 FILLER_46_1000 ();
 FILLCELL_X1 FILLER_46_1036 ();
 FILLCELL_X1 FILLER_46_1048 ();
 FILLCELL_X2 FILLER_46_1103 ();
 FILLCELL_X1 FILLER_46_1114 ();
 FILLCELL_X1 FILLER_47_33 ();
 FILLCELL_X4 FILLER_47_50 ();
 FILLCELL_X2 FILLER_47_54 ();
 FILLCELL_X1 FILLER_47_56 ();
 FILLCELL_X1 FILLER_47_71 ();
 FILLCELL_X4 FILLER_47_90 ();
 FILLCELL_X2 FILLER_47_94 ();
 FILLCELL_X1 FILLER_47_96 ();
 FILLCELL_X8 FILLER_47_115 ();
 FILLCELL_X2 FILLER_47_123 ();
 FILLCELL_X1 FILLER_47_125 ();
 FILLCELL_X1 FILLER_47_148 ();
 FILLCELL_X4 FILLER_47_153 ();
 FILLCELL_X2 FILLER_47_209 ();
 FILLCELL_X1 FILLER_47_211 ();
 FILLCELL_X1 FILLER_47_226 ();
 FILLCELL_X2 FILLER_47_241 ();
 FILLCELL_X1 FILLER_47_245 ();
 FILLCELL_X4 FILLER_47_262 ();
 FILLCELL_X2 FILLER_47_270 ();
 FILLCELL_X4 FILLER_47_294 ();
 FILLCELL_X1 FILLER_47_305 ();
 FILLCELL_X8 FILLER_47_360 ();
 FILLCELL_X1 FILLER_47_396 ();
 FILLCELL_X1 FILLER_47_546 ();
 FILLCELL_X1 FILLER_47_579 ();
 FILLCELL_X2 FILLER_47_626 ();
 FILLCELL_X1 FILLER_47_628 ();
 FILLCELL_X8 FILLER_47_649 ();
 FILLCELL_X4 FILLER_47_657 ();
 FILLCELL_X1 FILLER_47_661 ();
 FILLCELL_X4 FILLER_47_676 ();
 FILLCELL_X2 FILLER_47_680 ();
 FILLCELL_X1 FILLER_47_682 ();
 FILLCELL_X4 FILLER_47_687 ();
 FILLCELL_X2 FILLER_47_695 ();
 FILLCELL_X2 FILLER_47_701 ();
 FILLCELL_X1 FILLER_47_709 ();
 FILLCELL_X2 FILLER_47_725 ();
 FILLCELL_X1 FILLER_47_727 ();
 FILLCELL_X8 FILLER_47_768 ();
 FILLCELL_X2 FILLER_47_798 ();
 FILLCELL_X16 FILLER_47_802 ();
 FILLCELL_X2 FILLER_47_828 ();
 FILLCELL_X2 FILLER_47_845 ();
 FILLCELL_X1 FILLER_47_847 ();
 FILLCELL_X1 FILLER_47_913 ();
 FILLCELL_X1 FILLER_47_934 ();
 FILLCELL_X1 FILLER_47_940 ();
 FILLCELL_X1 FILLER_47_947 ();
 FILLCELL_X1 FILLER_47_955 ();
 FILLCELL_X1 FILLER_47_965 ();
 FILLCELL_X1 FILLER_47_968 ();
 FILLCELL_X2 FILLER_47_979 ();
 FILLCELL_X2 FILLER_47_986 ();
 FILLCELL_X1 FILLER_47_988 ();
 FILLCELL_X1 FILLER_47_998 ();
 FILLCELL_X1 FILLER_47_1033 ();
 FILLCELL_X2 FILLER_47_1038 ();
 FILLCELL_X2 FILLER_47_1043 ();
 FILLCELL_X2 FILLER_47_1049 ();
 FILLCELL_X1 FILLER_47_1057 ();
 FILLCELL_X1 FILLER_47_1083 ();
 FILLCELL_X1 FILLER_47_1098 ();
 FILLCELL_X1 FILLER_47_1115 ();
 FILLCELL_X1 FILLER_48_21 ();
 FILLCELL_X1 FILLER_48_56 ();
 FILLCELL_X1 FILLER_48_73 ();
 FILLCELL_X4 FILLER_48_100 ();
 FILLCELL_X2 FILLER_48_104 ();
 FILLCELL_X4 FILLER_48_114 ();
 FILLCELL_X2 FILLER_48_118 ();
 FILLCELL_X2 FILLER_48_123 ();
 FILLCELL_X1 FILLER_48_125 ();
 FILLCELL_X4 FILLER_48_133 ();
 FILLCELL_X2 FILLER_48_137 ();
 FILLCELL_X1 FILLER_48_163 ();
 FILLCELL_X2 FILLER_48_170 ();
 FILLCELL_X1 FILLER_48_172 ();
 FILLCELL_X8 FILLER_48_189 ();
 FILLCELL_X1 FILLER_48_197 ();
 FILLCELL_X32 FILLER_48_268 ();
 FILLCELL_X2 FILLER_48_300 ();
 FILLCELL_X1 FILLER_48_302 ();
 FILLCELL_X1 FILLER_48_311 ();
 FILLCELL_X1 FILLER_48_385 ();
 FILLCELL_X2 FILLER_48_393 ();
 FILLCELL_X2 FILLER_48_619 ();
 FILLCELL_X2 FILLER_48_642 ();
 FILLCELL_X1 FILLER_48_644 ();
 FILLCELL_X1 FILLER_48_659 ();
 FILLCELL_X2 FILLER_48_664 ();
 FILLCELL_X1 FILLER_48_697 ();
 FILLCELL_X2 FILLER_48_723 ();
 FILLCELL_X2 FILLER_48_745 ();
 FILLCELL_X1 FILLER_48_747 ();
 FILLCELL_X2 FILLER_48_819 ();
 FILLCELL_X1 FILLER_48_823 ();
 FILLCELL_X1 FILLER_48_826 ();
 FILLCELL_X2 FILLER_48_831 ();
 FILLCELL_X4 FILLER_48_861 ();
 FILLCELL_X1 FILLER_48_897 ();
 FILLCELL_X1 FILLER_48_903 ();
 FILLCELL_X8 FILLER_48_917 ();
 FILLCELL_X2 FILLER_48_925 ();
 FILLCELL_X4 FILLER_48_948 ();
 FILLCELL_X2 FILLER_48_952 ();
 FILLCELL_X1 FILLER_48_1030 ();
 FILLCELL_X4 FILLER_48_1035 ();
 FILLCELL_X1 FILLER_48_1061 ();
 FILLCELL_X2 FILLER_48_1139 ();
 FILLCELL_X2 FILLER_48_1146 ();
 FILLCELL_X2 FILLER_49_29 ();
 FILLCELL_X1 FILLER_49_35 ();
 FILLCELL_X8 FILLER_49_40 ();
 FILLCELL_X4 FILLER_49_48 ();
 FILLCELL_X2 FILLER_49_52 ();
 FILLCELL_X8 FILLER_49_58 ();
 FILLCELL_X1 FILLER_49_66 ();
 FILLCELL_X4 FILLER_49_79 ();
 FILLCELL_X2 FILLER_49_83 ();
 FILLCELL_X1 FILLER_49_85 ();
 FILLCELL_X1 FILLER_49_102 ();
 FILLCELL_X1 FILLER_49_135 ();
 FILLCELL_X1 FILLER_49_140 ();
 FILLCELL_X2 FILLER_49_151 ();
 FILLCELL_X1 FILLER_49_155 ();
 FILLCELL_X8 FILLER_49_172 ();
 FILLCELL_X4 FILLER_49_180 ();
 FILLCELL_X1 FILLER_49_184 ();
 FILLCELL_X8 FILLER_49_187 ();
 FILLCELL_X4 FILLER_49_195 ();
 FILLCELL_X8 FILLER_49_222 ();
 FILLCELL_X1 FILLER_49_230 ();
 FILLCELL_X4 FILLER_49_233 ();
 FILLCELL_X4 FILLER_49_249 ();
 FILLCELL_X1 FILLER_49_253 ();
 FILLCELL_X4 FILLER_49_256 ();
 FILLCELL_X2 FILLER_49_260 ();
 FILLCELL_X1 FILLER_49_262 ();
 FILLCELL_X2 FILLER_49_265 ();
 FILLCELL_X1 FILLER_49_267 ();
 FILLCELL_X4 FILLER_49_270 ();
 FILLCELL_X2 FILLER_49_274 ();
 FILLCELL_X2 FILLER_49_296 ();
 FILLCELL_X1 FILLER_49_310 ();
 FILLCELL_X1 FILLER_49_333 ();
 FILLCELL_X2 FILLER_49_337 ();
 FILLCELL_X2 FILLER_49_378 ();
 FILLCELL_X1 FILLER_49_422 ();
 FILLCELL_X1 FILLER_49_435 ();
 FILLCELL_X1 FILLER_49_569 ();
 FILLCELL_X1 FILLER_49_616 ();
 FILLCELL_X1 FILLER_49_627 ();
 FILLCELL_X1 FILLER_49_634 ();
 FILLCELL_X2 FILLER_49_639 ();
 FILLCELL_X2 FILLER_49_644 ();
 FILLCELL_X2 FILLER_49_650 ();
 FILLCELL_X2 FILLER_49_670 ();
 FILLCELL_X1 FILLER_49_714 ();
 FILLCELL_X2 FILLER_49_733 ();
 FILLCELL_X4 FILLER_49_745 ();
 FILLCELL_X1 FILLER_49_749 ();
 FILLCELL_X4 FILLER_49_766 ();
 FILLCELL_X1 FILLER_49_770 ();
 FILLCELL_X1 FILLER_49_773 ();
 FILLCELL_X1 FILLER_49_794 ();
 FILLCELL_X2 FILLER_49_805 ();
 FILLCELL_X4 FILLER_49_815 ();
 FILLCELL_X2 FILLER_49_829 ();
 FILLCELL_X2 FILLER_49_862 ();
 FILLCELL_X1 FILLER_49_864 ();
 FILLCELL_X2 FILLER_49_893 ();
 FILLCELL_X2 FILLER_49_899 ();
 FILLCELL_X1 FILLER_49_931 ();
 FILLCELL_X4 FILLER_49_944 ();
 FILLCELL_X2 FILLER_49_948 ();
 FILLCELL_X2 FILLER_49_996 ();
 FILLCELL_X2 FILLER_49_1012 ();
 FILLCELL_X2 FILLER_49_1017 ();
 FILLCELL_X1 FILLER_49_1019 ();
 FILLCELL_X1 FILLER_49_1027 ();
 FILLCELL_X2 FILLER_49_1032 ();
 FILLCELL_X1 FILLER_49_1034 ();
 FILLCELL_X1 FILLER_49_1100 ();
 FILLCELL_X1 FILLER_49_1147 ();
 FILLCELL_X1 FILLER_50_4 ();
 FILLCELL_X1 FILLER_50_46 ();
 FILLCELL_X1 FILLER_50_63 ();
 FILLCELL_X1 FILLER_50_66 ();
 FILLCELL_X4 FILLER_50_83 ();
 FILLCELL_X2 FILLER_50_87 ();
 FILLCELL_X1 FILLER_50_89 ();
 FILLCELL_X1 FILLER_50_94 ();
 FILLCELL_X4 FILLER_50_101 ();
 FILLCELL_X2 FILLER_50_105 ();
 FILLCELL_X2 FILLER_50_115 ();
 FILLCELL_X1 FILLER_50_117 ();
 FILLCELL_X4 FILLER_50_120 ();
 FILLCELL_X1 FILLER_50_130 ();
 FILLCELL_X1 FILLER_50_162 ();
 FILLCELL_X2 FILLER_50_175 ();
 FILLCELL_X4 FILLER_50_212 ();
 FILLCELL_X1 FILLER_50_216 ();
 FILLCELL_X16 FILLER_50_253 ();
 FILLCELL_X4 FILLER_50_269 ();
 FILLCELL_X4 FILLER_50_293 ();
 FILLCELL_X2 FILLER_50_297 ();
 FILLCELL_X4 FILLER_50_335 ();
 FILLCELL_X4 FILLER_50_342 ();
 FILLCELL_X2 FILLER_50_346 ();
 FILLCELL_X1 FILLER_50_370 ();
 FILLCELL_X1 FILLER_50_385 ();
 FILLCELL_X1 FILLER_50_389 ();
 FILLCELL_X1 FILLER_50_422 ();
 FILLCELL_X2 FILLER_50_486 ();
 FILLCELL_X1 FILLER_50_578 ();
 FILLCELL_X2 FILLER_50_584 ();
 FILLCELL_X4 FILLER_50_602 ();
 FILLCELL_X8 FILLER_50_608 ();
 FILLCELL_X4 FILLER_50_616 ();
 FILLCELL_X4 FILLER_50_624 ();
 FILLCELL_X1 FILLER_50_628 ();
 FILLCELL_X2 FILLER_50_662 ();
 FILLCELL_X1 FILLER_50_664 ();
 FILLCELL_X2 FILLER_50_687 ();
 FILLCELL_X1 FILLER_50_689 ();
 FILLCELL_X1 FILLER_50_725 ();
 FILLCELL_X1 FILLER_50_740 ();
 FILLCELL_X2 FILLER_50_767 ();
 FILLCELL_X1 FILLER_50_769 ();
 FILLCELL_X4 FILLER_50_790 ();
 FILLCELL_X2 FILLER_50_794 ();
 FILLCELL_X2 FILLER_50_806 ();
 FILLCELL_X1 FILLER_50_814 ();
 FILLCELL_X1 FILLER_50_887 ();
 FILLCELL_X1 FILLER_50_891 ();
 FILLCELL_X1 FILLER_50_894 ();
 FILLCELL_X4 FILLER_50_905 ();
 FILLCELL_X1 FILLER_50_909 ();
 FILLCELL_X1 FILLER_50_930 ();
 FILLCELL_X4 FILLER_50_949 ();
 FILLCELL_X1 FILLER_50_953 ();
 FILLCELL_X1 FILLER_50_959 ();
 FILLCELL_X1 FILLER_50_962 ();
 FILLCELL_X1 FILLER_50_975 ();
 FILLCELL_X1 FILLER_50_1024 ();
 FILLCELL_X1 FILLER_50_1029 ();
 FILLCELL_X1 FILLER_50_1034 ();
 FILLCELL_X1 FILLER_50_1039 ();
 FILLCELL_X1 FILLER_50_1096 ();
 FILLCELL_X1 FILLER_50_1133 ();
 FILLCELL_X2 FILLER_51_17 ();
 FILLCELL_X1 FILLER_51_19 ();
 FILLCELL_X8 FILLER_51_59 ();
 FILLCELL_X4 FILLER_51_67 ();
 FILLCELL_X1 FILLER_51_110 ();
 FILLCELL_X1 FILLER_51_119 ();
 FILLCELL_X2 FILLER_51_138 ();
 FILLCELL_X2 FILLER_51_188 ();
 FILLCELL_X1 FILLER_51_190 ();
 FILLCELL_X2 FILLER_51_261 ();
 FILLCELL_X2 FILLER_51_290 ();
 FILLCELL_X1 FILLER_51_318 ();
 FILLCELL_X4 FILLER_51_333 ();
 FILLCELL_X2 FILLER_51_357 ();
 FILLCELL_X1 FILLER_51_396 ();
 FILLCELL_X1 FILLER_51_414 ();
 FILLCELL_X4 FILLER_51_422 ();
 FILLCELL_X2 FILLER_51_508 ();
 FILLCELL_X1 FILLER_51_510 ();
 FILLCELL_X1 FILLER_51_558 ();
 FILLCELL_X1 FILLER_51_580 ();
 FILLCELL_X2 FILLER_51_583 ();
 FILLCELL_X1 FILLER_51_601 ();
 FILLCELL_X2 FILLER_51_622 ();
 FILLCELL_X1 FILLER_51_624 ();
 FILLCELL_X2 FILLER_51_658 ();
 FILLCELL_X1 FILLER_51_683 ();
 FILLCELL_X1 FILLER_51_694 ();
 FILLCELL_X2 FILLER_51_699 ();
 FILLCELL_X2 FILLER_51_709 ();
 FILLCELL_X1 FILLER_51_722 ();
 FILLCELL_X2 FILLER_51_729 ();
 FILLCELL_X1 FILLER_51_739 ();
 FILLCELL_X4 FILLER_51_745 ();
 FILLCELL_X1 FILLER_51_749 ();
 FILLCELL_X2 FILLER_51_768 ();
 FILLCELL_X1 FILLER_51_770 ();
 FILLCELL_X1 FILLER_51_791 ();
 FILLCELL_X2 FILLER_51_802 ();
 FILLCELL_X1 FILLER_51_811 ();
 FILLCELL_X1 FILLER_51_834 ();
 FILLCELL_X2 FILLER_51_839 ();
 FILLCELL_X1 FILLER_51_841 ();
 FILLCELL_X4 FILLER_51_879 ();
 FILLCELL_X2 FILLER_51_886 ();
 FILLCELL_X1 FILLER_51_888 ();
 FILLCELL_X2 FILLER_51_913 ();
 FILLCELL_X4 FILLER_51_925 ();
 FILLCELL_X2 FILLER_51_929 ();
 FILLCELL_X1 FILLER_51_931 ();
 FILLCELL_X1 FILLER_51_936 ();
 FILLCELL_X1 FILLER_51_939 ();
 FILLCELL_X4 FILLER_51_950 ();
 FILLCELL_X1 FILLER_51_954 ();
 FILLCELL_X1 FILLER_51_1012 ();
 FILLCELL_X1 FILLER_51_1022 ();
 FILLCELL_X1 FILLER_51_1026 ();
 FILLCELL_X1 FILLER_51_1049 ();
 FILLCELL_X1 FILLER_51_1070 ();
 FILLCELL_X1 FILLER_51_1089 ();
 FILLCELL_X1 FILLER_52_22 ();
 FILLCELL_X2 FILLER_52_26 ();
 FILLCELL_X1 FILLER_52_44 ();
 FILLCELL_X4 FILLER_52_47 ();
 FILLCELL_X2 FILLER_52_53 ();
 FILLCELL_X2 FILLER_52_57 ();
 FILLCELL_X2 FILLER_52_67 ();
 FILLCELL_X2 FILLER_52_85 ();
 FILLCELL_X1 FILLER_52_105 ();
 FILLCELL_X2 FILLER_52_122 ();
 FILLCELL_X1 FILLER_52_124 ();
 FILLCELL_X2 FILLER_52_130 ();
 FILLCELL_X1 FILLER_52_136 ();
 FILLCELL_X2 FILLER_52_141 ();
 FILLCELL_X2 FILLER_52_147 ();
 FILLCELL_X1 FILLER_52_153 ();
 FILLCELL_X2 FILLER_52_193 ();
 FILLCELL_X8 FILLER_52_199 ();
 FILLCELL_X2 FILLER_52_207 ();
 FILLCELL_X1 FILLER_52_211 ();
 FILLCELL_X1 FILLER_52_228 ();
 FILLCELL_X1 FILLER_52_245 ();
 FILLCELL_X1 FILLER_52_326 ();
 FILLCELL_X2 FILLER_52_334 ();
 FILLCELL_X2 FILLER_52_368 ();
 FILLCELL_X1 FILLER_52_370 ();
 FILLCELL_X2 FILLER_52_404 ();
 FILLCELL_X1 FILLER_52_413 ();
 FILLCELL_X1 FILLER_52_572 ();
 FILLCELL_X8 FILLER_52_579 ();
 FILLCELL_X2 FILLER_52_587 ();
 FILLCELL_X2 FILLER_52_611 ();
 FILLCELL_X4 FILLER_52_623 ();
 FILLCELL_X1 FILLER_52_641 ();
 FILLCELL_X1 FILLER_52_645 ();
 FILLCELL_X4 FILLER_52_663 ();
 FILLCELL_X1 FILLER_52_689 ();
 FILLCELL_X16 FILLER_52_702 ();
 FILLCELL_X4 FILLER_52_744 ();
 FILLCELL_X2 FILLER_52_748 ();
 FILLCELL_X1 FILLER_52_821 ();
 FILLCELL_X1 FILLER_52_841 ();
 FILLCELL_X1 FILLER_52_880 ();
 FILLCELL_X1 FILLER_52_912 ();
 FILLCELL_X2 FILLER_52_936 ();
 FILLCELL_X1 FILLER_52_951 ();
 FILLCELL_X1 FILLER_52_956 ();
 FILLCELL_X2 FILLER_52_990 ();
 FILLCELL_X1 FILLER_52_1123 ();
 FILLCELL_X1 FILLER_52_1142 ();
 FILLCELL_X4 FILLER_53_1 ();
 FILLCELL_X2 FILLER_53_5 ();
 FILLCELL_X1 FILLER_53_7 ();
 FILLCELL_X4 FILLER_53_15 ();
 FILLCELL_X2 FILLER_53_19 ();
 FILLCELL_X1 FILLER_53_21 ();
 FILLCELL_X4 FILLER_53_31 ();
 FILLCELL_X2 FILLER_53_85 ();
 FILLCELL_X1 FILLER_53_87 ();
 FILLCELL_X2 FILLER_53_90 ();
 FILLCELL_X1 FILLER_53_92 ();
 FILLCELL_X1 FILLER_53_143 ();
 FILLCELL_X1 FILLER_53_148 ();
 FILLCELL_X2 FILLER_53_159 ();
 FILLCELL_X1 FILLER_53_161 ();
 FILLCELL_X1 FILLER_53_180 ();
 FILLCELL_X8 FILLER_53_203 ();
 FILLCELL_X2 FILLER_53_211 ();
 FILLCELL_X1 FILLER_53_213 ();
 FILLCELL_X1 FILLER_53_216 ();
 FILLCELL_X4 FILLER_53_235 ();
 FILLCELL_X2 FILLER_53_259 ();
 FILLCELL_X1 FILLER_53_293 ();
 FILLCELL_X1 FILLER_53_298 ();
 FILLCELL_X1 FILLER_53_306 ();
 FILLCELL_X1 FILLER_53_309 ();
 FILLCELL_X1 FILLER_53_336 ();
 FILLCELL_X1 FILLER_53_340 ();
 FILLCELL_X8 FILLER_53_349 ();
 FILLCELL_X4 FILLER_53_357 ();
 FILLCELL_X2 FILLER_53_361 ();
 FILLCELL_X1 FILLER_53_363 ();
 FILLCELL_X1 FILLER_53_382 ();
 FILLCELL_X1 FILLER_53_390 ();
 FILLCELL_X1 FILLER_53_402 ();
 FILLCELL_X1 FILLER_53_413 ();
 FILLCELL_X1 FILLER_53_520 ();
 FILLCELL_X2 FILLER_53_556 ();
 FILLCELL_X1 FILLER_53_558 ();
 FILLCELL_X1 FILLER_53_581 ();
 FILLCELL_X4 FILLER_53_585 ();
 FILLCELL_X2 FILLER_53_589 ();
 FILLCELL_X1 FILLER_53_613 ();
 FILLCELL_X2 FILLER_53_618 ();
 FILLCELL_X1 FILLER_53_620 ();
 FILLCELL_X2 FILLER_53_624 ();
 FILLCELL_X1 FILLER_53_626 ();
 FILLCELL_X2 FILLER_53_647 ();
 FILLCELL_X2 FILLER_53_656 ();
 FILLCELL_X2 FILLER_53_669 ();
 FILLCELL_X4 FILLER_53_688 ();
 FILLCELL_X1 FILLER_53_714 ();
 FILLCELL_X1 FILLER_53_745 ();
 FILLCELL_X16 FILLER_53_753 ();
 FILLCELL_X2 FILLER_53_771 ();
 FILLCELL_X8 FILLER_53_776 ();
 FILLCELL_X4 FILLER_53_784 ();
 FILLCELL_X1 FILLER_53_788 ();
 FILLCELL_X4 FILLER_53_821 ();
 FILLCELL_X1 FILLER_53_825 ();
 FILLCELL_X1 FILLER_53_830 ();
 FILLCELL_X1 FILLER_53_843 ();
 FILLCELL_X2 FILLER_53_850 ();
 FILLCELL_X1 FILLER_53_852 ();
 FILLCELL_X1 FILLER_53_867 ();
 FILLCELL_X1 FILLER_53_888 ();
 FILLCELL_X1 FILLER_53_899 ();
 FILLCELL_X1 FILLER_53_903 ();
 FILLCELL_X2 FILLER_53_911 ();
 FILLCELL_X1 FILLER_53_933 ();
 FILLCELL_X2 FILLER_53_947 ();
 FILLCELL_X1 FILLER_53_949 ();
 FILLCELL_X1 FILLER_53_1076 ();
 FILLCELL_X1 FILLER_53_1084 ();
 FILLCELL_X1 FILLER_53_1128 ();
 FILLCELL_X1 FILLER_54_1 ();
 FILLCELL_X8 FILLER_54_5 ();
 FILLCELL_X1 FILLER_54_13 ();
 FILLCELL_X8 FILLER_54_30 ();
 FILLCELL_X4 FILLER_54_38 ();
 FILLCELL_X1 FILLER_54_70 ();
 FILLCELL_X4 FILLER_54_73 ();
 FILLCELL_X2 FILLER_54_77 ();
 FILLCELL_X1 FILLER_54_79 ();
 FILLCELL_X8 FILLER_54_96 ();
 FILLCELL_X4 FILLER_54_108 ();
 FILLCELL_X2 FILLER_54_112 ();
 FILLCELL_X2 FILLER_54_133 ();
 FILLCELL_X2 FILLER_54_143 ();
 FILLCELL_X1 FILLER_54_145 ();
 FILLCELL_X4 FILLER_54_154 ();
 FILLCELL_X2 FILLER_54_158 ();
 FILLCELL_X2 FILLER_54_164 ();
 FILLCELL_X2 FILLER_54_192 ();
 FILLCELL_X1 FILLER_54_194 ();
 FILLCELL_X4 FILLER_54_198 ();
 FILLCELL_X4 FILLER_54_222 ();
 FILLCELL_X4 FILLER_54_228 ();
 FILLCELL_X2 FILLER_54_232 ();
 FILLCELL_X2 FILLER_54_276 ();
 FILLCELL_X1 FILLER_54_278 ();
 FILLCELL_X1 FILLER_54_297 ();
 FILLCELL_X1 FILLER_54_302 ();
 FILLCELL_X1 FILLER_54_315 ();
 FILLCELL_X1 FILLER_54_386 ();
 FILLCELL_X1 FILLER_54_389 ();
 FILLCELL_X1 FILLER_54_401 ();
 FILLCELL_X2 FILLER_54_504 ();
 FILLCELL_X1 FILLER_54_542 ();
 FILLCELL_X1 FILLER_54_589 ();
 FILLCELL_X1 FILLER_54_610 ();
 FILLCELL_X1 FILLER_54_668 ();
 FILLCELL_X1 FILLER_54_688 ();
 FILLCELL_X4 FILLER_54_699 ();
 FILLCELL_X1 FILLER_54_728 ();
 FILLCELL_X4 FILLER_54_745 ();
 FILLCELL_X2 FILLER_54_759 ();
 FILLCELL_X1 FILLER_54_813 ();
 FILLCELL_X2 FILLER_54_833 ();
 FILLCELL_X1 FILLER_54_849 ();
 FILLCELL_X1 FILLER_54_860 ();
 FILLCELL_X1 FILLER_54_899 ();
 FILLCELL_X1 FILLER_54_948 ();
 FILLCELL_X1 FILLER_54_981 ();
 FILLCELL_X2 FILLER_54_1022 ();
 FILLCELL_X1 FILLER_54_1049 ();
 FILLCELL_X1 FILLER_54_1074 ();
 FILLCELL_X2 FILLER_54_1136 ();
 FILLCELL_X1 FILLER_54_1138 ();
 FILLCELL_X8 FILLER_55_5 ();
 FILLCELL_X4 FILLER_55_13 ();
 FILLCELL_X8 FILLER_55_21 ();
 FILLCELL_X1 FILLER_55_47 ();
 FILLCELL_X8 FILLER_55_112 ();
 FILLCELL_X4 FILLER_55_120 ();
 FILLCELL_X1 FILLER_55_158 ();
 FILLCELL_X1 FILLER_55_171 ();
 FILLCELL_X2 FILLER_55_180 ();
 FILLCELL_X1 FILLER_55_186 ();
 FILLCELL_X2 FILLER_55_205 ();
 FILLCELL_X16 FILLER_55_209 ();
 FILLCELL_X8 FILLER_55_225 ();
 FILLCELL_X4 FILLER_55_253 ();
 FILLCELL_X2 FILLER_55_257 ();
 FILLCELL_X1 FILLER_55_259 ();
 FILLCELL_X1 FILLER_55_298 ();
 FILLCELL_X2 FILLER_55_314 ();
 FILLCELL_X1 FILLER_55_316 ();
 FILLCELL_X1 FILLER_55_321 ();
 FILLCELL_X2 FILLER_55_333 ();
 FILLCELL_X2 FILLER_55_358 ();
 FILLCELL_X2 FILLER_55_409 ();
 FILLCELL_X1 FILLER_55_488 ();
 FILLCELL_X1 FILLER_55_532 ();
 FILLCELL_X2 FILLER_55_571 ();
 FILLCELL_X1 FILLER_55_577 ();
 FILLCELL_X4 FILLER_55_582 ();
 FILLCELL_X1 FILLER_55_586 ();
 FILLCELL_X1 FILLER_55_628 ();
 FILLCELL_X1 FILLER_55_633 ();
 FILLCELL_X1 FILLER_55_641 ();
 FILLCELL_X1 FILLER_55_674 ();
 FILLCELL_X1 FILLER_55_685 ();
 FILLCELL_X4 FILLER_55_696 ();
 FILLCELL_X4 FILLER_55_729 ();
 FILLCELL_X1 FILLER_55_733 ();
 FILLCELL_X1 FILLER_55_840 ();
 FILLCELL_X1 FILLER_55_874 ();
 FILLCELL_X1 FILLER_55_898 ();
 FILLCELL_X1 FILLER_55_902 ();
 FILLCELL_X1 FILLER_55_906 ();
 FILLCELL_X2 FILLER_55_1048 ();
 FILLCELL_X2 FILLER_55_1138 ();
 FILLCELL_X1 FILLER_55_1140 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X8 FILLER_56_35 ();
 FILLCELL_X2 FILLER_56_43 ();
 FILLCELL_X1 FILLER_56_45 ();
 FILLCELL_X4 FILLER_56_50 ();
 FILLCELL_X1 FILLER_56_54 ();
 FILLCELL_X4 FILLER_56_58 ();
 FILLCELL_X2 FILLER_56_62 ();
 FILLCELL_X1 FILLER_56_146 ();
 FILLCELL_X4 FILLER_56_163 ();
 FILLCELL_X2 FILLER_56_183 ();
 FILLCELL_X1 FILLER_56_189 ();
 FILLCELL_X4 FILLER_56_210 ();
 FILLCELL_X4 FILLER_56_236 ();
 FILLCELL_X2 FILLER_56_240 ();
 FILLCELL_X1 FILLER_56_247 ();
 FILLCELL_X4 FILLER_56_268 ();
 FILLCELL_X2 FILLER_56_272 ();
 FILLCELL_X1 FILLER_56_288 ();
 FILLCELL_X1 FILLER_56_311 ();
 FILLCELL_X4 FILLER_56_318 ();
 FILLCELL_X1 FILLER_56_359 ();
 FILLCELL_X1 FILLER_56_377 ();
 FILLCELL_X2 FILLER_56_395 ();
 FILLCELL_X2 FILLER_56_425 ();
 FILLCELL_X1 FILLER_56_427 ();
 FILLCELL_X2 FILLER_56_452 ();
 FILLCELL_X2 FILLER_56_497 ();
 FILLCELL_X1 FILLER_56_499 ();
 FILLCELL_X1 FILLER_56_503 ();
 FILLCELL_X2 FILLER_56_577 ();
 FILLCELL_X1 FILLER_56_579 ();
 FILLCELL_X4 FILLER_56_588 ();
 FILLCELL_X4 FILLER_56_602 ();
 FILLCELL_X2 FILLER_56_606 ();
 FILLCELL_X4 FILLER_56_612 ();
 FILLCELL_X2 FILLER_56_616 ();
 FILLCELL_X1 FILLER_56_618 ();
 FILLCELL_X2 FILLER_56_657 ();
 FILLCELL_X2 FILLER_56_671 ();
 FILLCELL_X1 FILLER_56_673 ();
 FILLCELL_X2 FILLER_56_681 ();
 FILLCELL_X8 FILLER_56_709 ();
 FILLCELL_X8 FILLER_56_719 ();
 FILLCELL_X4 FILLER_56_727 ();
 FILLCELL_X2 FILLER_56_745 ();
 FILLCELL_X1 FILLER_56_747 ();
 FILLCELL_X1 FILLER_56_755 ();
 FILLCELL_X1 FILLER_56_783 ();
 FILLCELL_X1 FILLER_56_808 ();
 FILLCELL_X1 FILLER_56_903 ();
 FILLCELL_X2 FILLER_56_927 ();
 FILLCELL_X2 FILLER_56_963 ();
 FILLCELL_X1 FILLER_56_1002 ();
 FILLCELL_X1 FILLER_56_1027 ();
 FILLCELL_X1 FILLER_56_1044 ();
 FILLCELL_X1 FILLER_56_1063 ();
 FILLCELL_X1 FILLER_56_1075 ();
 FILLCELL_X1 FILLER_56_1085 ();
 FILLCELL_X1 FILLER_56_1093 ();
 FILLCELL_X1 FILLER_56_1117 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X8 FILLER_57_33 ();
 FILLCELL_X4 FILLER_57_41 ();
 FILLCELL_X1 FILLER_57_45 ();
 FILLCELL_X1 FILLER_57_62 ();
 FILLCELL_X2 FILLER_57_83 ();
 FILLCELL_X4 FILLER_57_87 ();
 FILLCELL_X2 FILLER_57_133 ();
 FILLCELL_X8 FILLER_57_155 ();
 FILLCELL_X16 FILLER_57_165 ();
 FILLCELL_X4 FILLER_57_181 ();
 FILLCELL_X1 FILLER_57_185 ();
 FILLCELL_X4 FILLER_57_202 ();
 FILLCELL_X8 FILLER_57_210 ();
 FILLCELL_X2 FILLER_57_218 ();
 FILLCELL_X8 FILLER_57_244 ();
 FILLCELL_X1 FILLER_57_252 ();
 FILLCELL_X4 FILLER_57_273 ();
 FILLCELL_X2 FILLER_57_287 ();
 FILLCELL_X2 FILLER_57_300 ();
 FILLCELL_X2 FILLER_57_316 ();
 FILLCELL_X1 FILLER_57_335 ();
 FILLCELL_X2 FILLER_57_339 ();
 FILLCELL_X2 FILLER_57_361 ();
 FILLCELL_X2 FILLER_57_402 ();
 FILLCELL_X2 FILLER_57_416 ();
 FILLCELL_X1 FILLER_57_427 ();
 FILLCELL_X1 FILLER_57_441 ();
 FILLCELL_X1 FILLER_57_504 ();
 FILLCELL_X1 FILLER_57_515 ();
 FILLCELL_X2 FILLER_57_539 ();
 FILLCELL_X2 FILLER_57_546 ();
 FILLCELL_X2 FILLER_57_557 ();
 FILLCELL_X2 FILLER_57_570 ();
 FILLCELL_X1 FILLER_57_572 ();
 FILLCELL_X4 FILLER_57_586 ();
 FILLCELL_X2 FILLER_57_590 ();
 FILLCELL_X4 FILLER_57_612 ();
 FILLCELL_X2 FILLER_57_616 ();
 FILLCELL_X4 FILLER_57_676 ();
 FILLCELL_X2 FILLER_57_710 ();
 FILLCELL_X1 FILLER_57_712 ();
 FILLCELL_X4 FILLER_57_723 ();
 FILLCELL_X1 FILLER_57_727 ();
 FILLCELL_X2 FILLER_57_747 ();
 FILLCELL_X1 FILLER_57_857 ();
 FILLCELL_X1 FILLER_57_862 ();
 FILLCELL_X1 FILLER_57_866 ();
 FILLCELL_X1 FILLER_57_883 ();
 FILLCELL_X1 FILLER_57_891 ();
 FILLCELL_X1 FILLER_57_897 ();
 FILLCELL_X1 FILLER_57_905 ();
 FILLCELL_X2 FILLER_57_910 ();
 FILLCELL_X2 FILLER_57_934 ();
 FILLCELL_X2 FILLER_57_953 ();
 FILLCELL_X1 FILLER_57_955 ();
 FILLCELL_X1 FILLER_57_976 ();
 FILLCELL_X1 FILLER_57_980 ();
 FILLCELL_X1 FILLER_57_985 ();
 FILLCELL_X1 FILLER_57_1033 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X16 FILLER_58_33 ();
 FILLCELL_X2 FILLER_58_49 ();
 FILLCELL_X2 FILLER_58_53 ();
 FILLCELL_X4 FILLER_58_57 ();
 FILLCELL_X2 FILLER_58_61 ();
 FILLCELL_X1 FILLER_58_63 ();
 FILLCELL_X4 FILLER_58_66 ();
 FILLCELL_X2 FILLER_58_70 ();
 FILLCELL_X1 FILLER_58_134 ();
 FILLCELL_X8 FILLER_58_137 ();
 FILLCELL_X4 FILLER_58_145 ();
 FILLCELL_X2 FILLER_58_151 ();
 FILLCELL_X1 FILLER_58_153 ();
 FILLCELL_X1 FILLER_58_172 ();
 FILLCELL_X4 FILLER_58_189 ();
 FILLCELL_X2 FILLER_58_193 ();
 FILLCELL_X1 FILLER_58_195 ();
 FILLCELL_X8 FILLER_58_200 ();
 FILLCELL_X4 FILLER_58_224 ();
 FILLCELL_X1 FILLER_58_228 ();
 FILLCELL_X4 FILLER_58_233 ();
 FILLCELL_X2 FILLER_58_237 ();
 FILLCELL_X1 FILLER_58_239 ();
 FILLCELL_X2 FILLER_58_260 ();
 FILLCELL_X8 FILLER_58_264 ();
 FILLCELL_X2 FILLER_58_272 ();
 FILLCELL_X1 FILLER_58_274 ();
 FILLCELL_X1 FILLER_58_297 ();
 FILLCELL_X1 FILLER_58_328 ();
 FILLCELL_X1 FILLER_58_331 ();
 FILLCELL_X2 FILLER_58_342 ();
 FILLCELL_X8 FILLER_58_364 ();
 FILLCELL_X4 FILLER_58_372 ();
 FILLCELL_X1 FILLER_58_376 ();
 FILLCELL_X4 FILLER_58_398 ();
 FILLCELL_X2 FILLER_58_402 ();
 FILLCELL_X2 FILLER_58_406 ();
 FILLCELL_X1 FILLER_58_429 ();
 FILLCELL_X2 FILLER_58_461 ();
 FILLCELL_X2 FILLER_58_550 ();
 FILLCELL_X2 FILLER_58_576 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X1 FILLER_58_636 ();
 FILLCELL_X2 FILLER_58_657 ();
 FILLCELL_X1 FILLER_58_662 ();
 FILLCELL_X1 FILLER_58_670 ();
 FILLCELL_X1 FILLER_58_693 ();
 FILLCELL_X1 FILLER_58_708 ();
 FILLCELL_X4 FILLER_58_729 ();
 FILLCELL_X2 FILLER_58_733 ();
 FILLCELL_X2 FILLER_58_757 ();
 FILLCELL_X1 FILLER_58_759 ();
 FILLCELL_X1 FILLER_58_782 ();
 FILLCELL_X2 FILLER_58_836 ();
 FILLCELL_X1 FILLER_58_896 ();
 FILLCELL_X1 FILLER_58_901 ();
 FILLCELL_X1 FILLER_58_936 ();
 FILLCELL_X1 FILLER_58_947 ();
 FILLCELL_X4 FILLER_58_958 ();
 FILLCELL_X2 FILLER_58_962 ();
 FILLCELL_X8 FILLER_58_971 ();
 FILLCELL_X1 FILLER_58_987 ();
 FILLCELL_X2 FILLER_58_1028 ();
 FILLCELL_X2 FILLER_58_1096 ();
 FILLCELL_X1 FILLER_58_1117 ();
 FILLCELL_X2 FILLER_58_1121 ();
 FILLCELL_X4 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X8 FILLER_59_33 ();
 FILLCELL_X1 FILLER_59_41 ();
 FILLCELL_X8 FILLER_59_44 ();
 FILLCELL_X2 FILLER_59_52 ();
 FILLCELL_X1 FILLER_59_74 ();
 FILLCELL_X32 FILLER_59_78 ();
 FILLCELL_X16 FILLER_59_110 ();
 FILLCELL_X2 FILLER_59_126 ();
 FILLCELL_X2 FILLER_59_204 ();
 FILLCELL_X1 FILLER_59_206 ();
 FILLCELL_X4 FILLER_59_237 ();
 FILLCELL_X2 FILLER_59_241 ();
 FILLCELL_X2 FILLER_59_283 ();
 FILLCELL_X1 FILLER_59_285 ();
 FILLCELL_X4 FILLER_59_335 ();
 FILLCELL_X16 FILLER_59_344 ();
 FILLCELL_X8 FILLER_59_360 ();
 FILLCELL_X4 FILLER_59_368 ();
 FILLCELL_X1 FILLER_59_372 ();
 FILLCELL_X4 FILLER_59_393 ();
 FILLCELL_X8 FILLER_59_399 ();
 FILLCELL_X4 FILLER_59_419 ();
 FILLCELL_X2 FILLER_59_438 ();
 FILLCELL_X1 FILLER_59_440 ();
 FILLCELL_X2 FILLER_59_485 ();
 FILLCELL_X2 FILLER_59_542 ();
 FILLCELL_X1 FILLER_59_544 ();
 FILLCELL_X4 FILLER_59_552 ();
 FILLCELL_X1 FILLER_59_556 ();
 FILLCELL_X4 FILLER_59_560 ();
 FILLCELL_X4 FILLER_59_570 ();
 FILLCELL_X2 FILLER_59_574 ();
 FILLCELL_X1 FILLER_59_576 ();
 FILLCELL_X2 FILLER_59_586 ();
 FILLCELL_X1 FILLER_59_588 ();
 FILLCELL_X4 FILLER_59_599 ();
 FILLCELL_X2 FILLER_59_649 ();
 FILLCELL_X1 FILLER_59_662 ();
 FILLCELL_X1 FILLER_59_670 ();
 FILLCELL_X1 FILLER_59_701 ();
 FILLCELL_X1 FILLER_59_712 ();
 FILLCELL_X8 FILLER_59_719 ();
 FILLCELL_X4 FILLER_59_727 ();
 FILLCELL_X2 FILLER_59_731 ();
 FILLCELL_X1 FILLER_59_835 ();
 FILLCELL_X1 FILLER_59_897 ();
 FILLCELL_X2 FILLER_59_918 ();
 FILLCELL_X2 FILLER_59_955 ();
 FILLCELL_X4 FILLER_59_964 ();
 FILLCELL_X2 FILLER_59_968 ();
 FILLCELL_X1 FILLER_59_994 ();
 FILLCELL_X2 FILLER_59_1043 ();
 FILLCELL_X1 FILLER_59_1045 ();
 FILLCELL_X1 FILLER_59_1053 ();
 FILLCELL_X2 FILLER_59_1116 ();
 FILLCELL_X1 FILLER_59_1140 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X8 FILLER_60_33 ();
 FILLCELL_X4 FILLER_60_41 ();
 FILLCELL_X2 FILLER_60_45 ();
 FILLCELL_X4 FILLER_60_73 ();
 FILLCELL_X2 FILLER_60_77 ();
 FILLCELL_X4 FILLER_60_81 ();
 FILLCELL_X1 FILLER_60_85 ();
 FILLCELL_X1 FILLER_60_113 ();
 FILLCELL_X16 FILLER_60_161 ();
 FILLCELL_X2 FILLER_60_177 ();
 FILLCELL_X1 FILLER_60_179 ();
 FILLCELL_X4 FILLER_60_280 ();
 FILLCELL_X2 FILLER_60_284 ();
 FILLCELL_X1 FILLER_60_286 ();
 FILLCELL_X1 FILLER_60_297 ();
 FILLCELL_X1 FILLER_60_309 ();
 FILLCELL_X1 FILLER_60_318 ();
 FILLCELL_X4 FILLER_60_338 ();
 FILLCELL_X1 FILLER_60_347 ();
 FILLCELL_X32 FILLER_60_352 ();
 FILLCELL_X16 FILLER_60_384 ();
 FILLCELL_X4 FILLER_60_400 ();
 FILLCELL_X2 FILLER_60_404 ();
 FILLCELL_X1 FILLER_60_418 ();
 FILLCELL_X1 FILLER_60_434 ();
 FILLCELL_X1 FILLER_60_529 ();
 FILLCELL_X2 FILLER_60_542 ();
 FILLCELL_X1 FILLER_60_544 ();
 FILLCELL_X1 FILLER_60_549 ();
 FILLCELL_X4 FILLER_60_609 ();
 FILLCELL_X1 FILLER_60_613 ();
 FILLCELL_X2 FILLER_60_663 ();
 FILLCELL_X1 FILLER_60_668 ();
 FILLCELL_X1 FILLER_60_675 ();
 FILLCELL_X2 FILLER_60_696 ();
 FILLCELL_X1 FILLER_60_698 ();
 FILLCELL_X2 FILLER_60_709 ();
 FILLCELL_X1 FILLER_60_711 ();
 FILLCELL_X2 FILLER_60_732 ();
 FILLCELL_X1 FILLER_60_734 ();
 FILLCELL_X1 FILLER_60_762 ();
 FILLCELL_X1 FILLER_60_807 ();
 FILLCELL_X1 FILLER_60_823 ();
 FILLCELL_X1 FILLER_60_828 ();
 FILLCELL_X1 FILLER_60_838 ();
 FILLCELL_X4 FILLER_60_921 ();
 FILLCELL_X2 FILLER_60_925 ();
 FILLCELL_X2 FILLER_60_947 ();
 FILLCELL_X4 FILLER_60_965 ();
 FILLCELL_X1 FILLER_60_969 ();
 FILLCELL_X2 FILLER_60_1143 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X8 FILLER_61_33 ();
 FILLCELL_X1 FILLER_61_41 ();
 FILLCELL_X1 FILLER_61_67 ();
 FILLCELL_X2 FILLER_61_110 ();
 FILLCELL_X8 FILLER_61_122 ();
 FILLCELL_X1 FILLER_61_199 ();
 FILLCELL_X2 FILLER_61_220 ();
 FILLCELL_X1 FILLER_61_222 ();
 FILLCELL_X8 FILLER_61_225 ();
 FILLCELL_X1 FILLER_61_233 ();
 FILLCELL_X2 FILLER_61_286 ();
 FILLCELL_X2 FILLER_61_302 ();
 FILLCELL_X1 FILLER_61_308 ();
 FILLCELL_X2 FILLER_61_342 ();
 FILLCELL_X1 FILLER_61_350 ();
 FILLCELL_X32 FILLER_61_374 ();
 FILLCELL_X4 FILLER_61_406 ();
 FILLCELL_X1 FILLER_61_410 ();
 FILLCELL_X1 FILLER_61_477 ();
 FILLCELL_X1 FILLER_61_483 ();
 FILLCELL_X4 FILLER_61_566 ();
 FILLCELL_X2 FILLER_61_570 ();
 FILLCELL_X1 FILLER_61_582 ();
 FILLCELL_X2 FILLER_61_621 ();
 FILLCELL_X1 FILLER_61_635 ();
 FILLCELL_X4 FILLER_61_656 ();
 FILLCELL_X2 FILLER_61_664 ();
 FILLCELL_X1 FILLER_61_666 ();
 FILLCELL_X16 FILLER_61_671 ();
 FILLCELL_X1 FILLER_61_715 ();
 FILLCELL_X2 FILLER_61_730 ();
 FILLCELL_X2 FILLER_61_840 ();
 FILLCELL_X1 FILLER_61_849 ();
 FILLCELL_X1 FILLER_61_908 ();
 FILLCELL_X2 FILLER_61_930 ();
 FILLCELL_X1 FILLER_61_966 ();
 FILLCELL_X1 FILLER_61_969 ();
 FILLCELL_X1 FILLER_61_980 ();
 FILLCELL_X1 FILLER_61_990 ();
 FILLCELL_X1 FILLER_61_996 ();
 FILLCELL_X1 FILLER_61_1147 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X8 FILLER_62_33 ();
 FILLCELL_X2 FILLER_62_41 ();
 FILLCELL_X1 FILLER_62_65 ();
 FILLCELL_X1 FILLER_62_86 ();
 FILLCELL_X2 FILLER_62_107 ();
 FILLCELL_X1 FILLER_62_119 ();
 FILLCELL_X2 FILLER_62_123 ();
 FILLCELL_X1 FILLER_62_125 ();
 FILLCELL_X1 FILLER_62_131 ();
 FILLCELL_X2 FILLER_62_140 ();
 FILLCELL_X1 FILLER_62_177 ();
 FILLCELL_X8 FILLER_62_208 ();
 FILLCELL_X2 FILLER_62_216 ();
 FILLCELL_X8 FILLER_62_282 ();
 FILLCELL_X8 FILLER_62_300 ();
 FILLCELL_X1 FILLER_62_308 ();
 FILLCELL_X4 FILLER_62_335 ();
 FILLCELL_X2 FILLER_62_354 ();
 FILLCELL_X32 FILLER_62_362 ();
 FILLCELL_X32 FILLER_62_394 ();
 FILLCELL_X1 FILLER_62_426 ();
 FILLCELL_X4 FILLER_62_430 ();
 FILLCELL_X4 FILLER_62_438 ();
 FILLCELL_X2 FILLER_62_450 ();
 FILLCELL_X1 FILLER_62_502 ();
 FILLCELL_X1 FILLER_62_563 ();
 FILLCELL_X1 FILLER_62_614 ();
 FILLCELL_X1 FILLER_62_619 ();
 FILLCELL_X2 FILLER_62_624 ();
 FILLCELL_X2 FILLER_62_628 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X2 FILLER_62_641 ();
 FILLCELL_X2 FILLER_62_648 ();
 FILLCELL_X8 FILLER_62_657 ();
 FILLCELL_X1 FILLER_62_665 ();
 FILLCELL_X1 FILLER_62_686 ();
 FILLCELL_X2 FILLER_62_738 ();
 FILLCELL_X1 FILLER_62_826 ();
 FILLCELL_X1 FILLER_62_913 ();
 FILLCELL_X2 FILLER_62_921 ();
 FILLCELL_X1 FILLER_62_926 ();
 FILLCELL_X2 FILLER_62_933 ();
 FILLCELL_X1 FILLER_62_935 ();
 FILLCELL_X1 FILLER_62_939 ();
 FILLCELL_X4 FILLER_62_960 ();
 FILLCELL_X1 FILLER_62_1101 ();
 FILLCELL_X1 FILLER_62_1147 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X8 FILLER_63_33 ();
 FILLCELL_X2 FILLER_63_41 ();
 FILLCELL_X1 FILLER_63_43 ();
 FILLCELL_X8 FILLER_63_64 ();
 FILLCELL_X1 FILLER_63_72 ();
 FILLCELL_X2 FILLER_63_83 ();
 FILLCELL_X2 FILLER_63_99 ();
 FILLCELL_X1 FILLER_63_101 ();
 FILLCELL_X2 FILLER_63_116 ();
 FILLCELL_X2 FILLER_63_122 ();
 FILLCELL_X1 FILLER_63_124 ();
 FILLCELL_X1 FILLER_63_127 ();
 FILLCELL_X2 FILLER_63_155 ();
 FILLCELL_X1 FILLER_63_181 ();
 FILLCELL_X2 FILLER_63_192 ();
 FILLCELL_X2 FILLER_63_198 ();
 FILLCELL_X2 FILLER_63_204 ();
 FILLCELL_X2 FILLER_63_210 ();
 FILLCELL_X4 FILLER_63_244 ();
 FILLCELL_X1 FILLER_63_248 ();
 FILLCELL_X4 FILLER_63_251 ();
 FILLCELL_X1 FILLER_63_255 ();
 FILLCELL_X16 FILLER_63_264 ();
 FILLCELL_X1 FILLER_63_280 ();
 FILLCELL_X16 FILLER_63_284 ();
 FILLCELL_X2 FILLER_63_300 ();
 FILLCELL_X1 FILLER_63_304 ();
 FILLCELL_X2 FILLER_63_329 ();
 FILLCELL_X2 FILLER_63_350 ();
 FILLCELL_X1 FILLER_63_352 ();
 FILLCELL_X4 FILLER_63_355 ();
 FILLCELL_X2 FILLER_63_359 ();
 FILLCELL_X2 FILLER_63_381 ();
 FILLCELL_X1 FILLER_63_383 ();
 FILLCELL_X32 FILLER_63_396 ();
 FILLCELL_X8 FILLER_63_428 ();
 FILLCELL_X4 FILLER_63_436 ();
 FILLCELL_X4 FILLER_63_447 ();
 FILLCELL_X16 FILLER_63_454 ();
 FILLCELL_X4 FILLER_63_470 ();
 FILLCELL_X1 FILLER_63_474 ();
 FILLCELL_X4 FILLER_63_589 ();
 FILLCELL_X2 FILLER_63_607 ();
 FILLCELL_X1 FILLER_63_609 ();
 FILLCELL_X1 FILLER_63_618 ();
 FILLCELL_X4 FILLER_63_645 ();
 FILLCELL_X16 FILLER_63_664 ();
 FILLCELL_X4 FILLER_63_680 ();
 FILLCELL_X2 FILLER_63_684 ();
 FILLCELL_X1 FILLER_63_690 ();
 FILLCELL_X2 FILLER_63_728 ();
 FILLCELL_X2 FILLER_63_740 ();
 FILLCELL_X1 FILLER_63_815 ();
 FILLCELL_X1 FILLER_63_870 ();
 FILLCELL_X2 FILLER_63_983 ();
 FILLCELL_X1 FILLER_63_985 ();
 FILLCELL_X2 FILLER_63_1094 ();
 FILLCELL_X1 FILLER_63_1143 ();
 FILLCELL_X1 FILLER_63_1147 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X16 FILLER_64_33 ();
 FILLCELL_X8 FILLER_64_49 ();
 FILLCELL_X2 FILLER_64_77 ();
 FILLCELL_X1 FILLER_64_79 ();
 FILLCELL_X2 FILLER_64_90 ();
 FILLCELL_X1 FILLER_64_92 ();
 FILLCELL_X4 FILLER_64_97 ();
 FILLCELL_X2 FILLER_64_157 ();
 FILLCELL_X1 FILLER_64_159 ();
 FILLCELL_X2 FILLER_64_197 ();
 FILLCELL_X1 FILLER_64_201 ();
 FILLCELL_X2 FILLER_64_209 ();
 FILLCELL_X2 FILLER_64_215 ();
 FILLCELL_X1 FILLER_64_221 ();
 FILLCELL_X4 FILLER_64_240 ();
 FILLCELL_X1 FILLER_64_244 ();
 FILLCELL_X4 FILLER_64_277 ();
 FILLCELL_X2 FILLER_64_301 ();
 FILLCELL_X2 FILLER_64_328 ();
 FILLCELL_X1 FILLER_64_330 ();
 FILLCELL_X1 FILLER_64_339 ();
 FILLCELL_X1 FILLER_64_350 ();
 FILLCELL_X4 FILLER_64_379 ();
 FILLCELL_X2 FILLER_64_383 ();
 FILLCELL_X1 FILLER_64_385 ();
 FILLCELL_X2 FILLER_64_393 ();
 FILLCELL_X32 FILLER_64_411 ();
 FILLCELL_X16 FILLER_64_443 ();
 FILLCELL_X8 FILLER_64_459 ();
 FILLCELL_X8 FILLER_64_469 ();
 FILLCELL_X1 FILLER_64_549 ();
 FILLCELL_X2 FILLER_64_606 ();
 FILLCELL_X1 FILLER_64_608 ();
 FILLCELL_X8 FILLER_64_616 ();
 FILLCELL_X1 FILLER_64_630 ();
 FILLCELL_X4 FILLER_64_638 ();
 FILLCELL_X32 FILLER_64_648 ();
 FILLCELL_X4 FILLER_64_680 ();
 FILLCELL_X1 FILLER_64_684 ();
 FILLCELL_X1 FILLER_64_694 ();
 FILLCELL_X1 FILLER_64_699 ();
 FILLCELL_X1 FILLER_64_735 ();
 FILLCELL_X1 FILLER_64_748 ();
 FILLCELL_X1 FILLER_64_752 ();
 FILLCELL_X1 FILLER_64_806 ();
 FILLCELL_X1 FILLER_64_899 ();
 FILLCELL_X4 FILLER_64_921 ();
 FILLCELL_X1 FILLER_64_1052 ();
 FILLCELL_X1 FILLER_64_1131 ();
 FILLCELL_X4 FILLER_64_1142 ();
 FILLCELL_X2 FILLER_64_1146 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X8 FILLER_65_33 ();
 FILLCELL_X4 FILLER_65_41 ();
 FILLCELL_X2 FILLER_65_45 ();
 FILLCELL_X1 FILLER_65_47 ();
 FILLCELL_X4 FILLER_65_50 ();
 FILLCELL_X2 FILLER_65_54 ();
 FILLCELL_X4 FILLER_65_76 ();
 FILLCELL_X1 FILLER_65_84 ();
 FILLCELL_X2 FILLER_65_89 ();
 FILLCELL_X2 FILLER_65_96 ();
 FILLCELL_X2 FILLER_65_102 ();
 FILLCELL_X1 FILLER_65_104 ();
 FILLCELL_X2 FILLER_65_138 ();
 FILLCELL_X2 FILLER_65_148 ();
 FILLCELL_X1 FILLER_65_150 ();
 FILLCELL_X2 FILLER_65_178 ();
 FILLCELL_X1 FILLER_65_188 ();
 FILLCELL_X4 FILLER_65_193 ();
 FILLCELL_X1 FILLER_65_197 ();
 FILLCELL_X4 FILLER_65_210 ();
 FILLCELL_X1 FILLER_65_214 ();
 FILLCELL_X4 FILLER_65_223 ();
 FILLCELL_X8 FILLER_65_233 ();
 FILLCELL_X4 FILLER_65_241 ();
 FILLCELL_X2 FILLER_65_245 ();
 FILLCELL_X4 FILLER_65_281 ();
 FILLCELL_X2 FILLER_65_288 ();
 FILLCELL_X1 FILLER_65_290 ();
 FILLCELL_X1 FILLER_65_311 ();
 FILLCELL_X2 FILLER_65_314 ();
 FILLCELL_X1 FILLER_65_316 ();
 FILLCELL_X1 FILLER_65_336 ();
 FILLCELL_X2 FILLER_65_357 ();
 FILLCELL_X1 FILLER_65_359 ();
 FILLCELL_X16 FILLER_65_364 ();
 FILLCELL_X4 FILLER_65_380 ();
 FILLCELL_X1 FILLER_65_384 ();
 FILLCELL_X32 FILLER_65_398 ();
 FILLCELL_X8 FILLER_65_430 ();
 FILLCELL_X16 FILLER_65_440 ();
 FILLCELL_X8 FILLER_65_456 ();
 FILLCELL_X4 FILLER_65_464 ();
 FILLCELL_X4 FILLER_65_470 ();
 FILLCELL_X1 FILLER_65_474 ();
 FILLCELL_X1 FILLER_65_504 ();
 FILLCELL_X8 FILLER_65_599 ();
 FILLCELL_X2 FILLER_65_607 ();
 FILLCELL_X4 FILLER_65_615 ();
 FILLCELL_X2 FILLER_65_619 ();
 FILLCELL_X1 FILLER_65_621 ();
 FILLCELL_X1 FILLER_65_652 ();
 FILLCELL_X4 FILLER_65_656 ();
 FILLCELL_X16 FILLER_65_664 ();
 FILLCELL_X2 FILLER_65_692 ();
 FILLCELL_X1 FILLER_65_704 ();
 FILLCELL_X1 FILLER_65_790 ();
 FILLCELL_X1 FILLER_65_926 ();
 FILLCELL_X2 FILLER_65_930 ();
 FILLCELL_X1 FILLER_65_959 ();
 FILLCELL_X1 FILLER_65_975 ();
 FILLCELL_X1 FILLER_65_983 ();
 FILLCELL_X2 FILLER_65_1111 ();
 FILLCELL_X1 FILLER_65_1116 ();
 FILLCELL_X1 FILLER_65_1121 ();
 FILLCELL_X16 FILLER_65_1129 ();
 FILLCELL_X2 FILLER_65_1145 ();
 FILLCELL_X1 FILLER_65_1147 ();
 FILLCELL_X2 FILLER_66_1 ();
 FILLCELL_X16 FILLER_66_6 ();
 FILLCELL_X4 FILLER_66_22 ();
 FILLCELL_X1 FILLER_66_26 ();
 FILLCELL_X1 FILLER_66_47 ();
 FILLCELL_X1 FILLER_66_124 ();
 FILLCELL_X1 FILLER_66_128 ();
 FILLCELL_X1 FILLER_66_141 ();
 FILLCELL_X4 FILLER_66_148 ();
 FILLCELL_X1 FILLER_66_171 ();
 FILLCELL_X4 FILLER_66_188 ();
 FILLCELL_X2 FILLER_66_208 ();
 FILLCELL_X1 FILLER_66_210 ();
 FILLCELL_X8 FILLER_66_241 ();
 FILLCELL_X4 FILLER_66_249 ();
 FILLCELL_X2 FILLER_66_253 ();
 FILLCELL_X1 FILLER_66_255 ();
 FILLCELL_X1 FILLER_66_263 ();
 FILLCELL_X1 FILLER_66_268 ();
 FILLCELL_X2 FILLER_66_275 ();
 FILLCELL_X1 FILLER_66_277 ();
 FILLCELL_X2 FILLER_66_290 ();
 FILLCELL_X2 FILLER_66_299 ();
 FILLCELL_X1 FILLER_66_301 ();
 FILLCELL_X2 FILLER_66_311 ();
 FILLCELL_X1 FILLER_66_313 ();
 FILLCELL_X2 FILLER_66_321 ();
 FILLCELL_X1 FILLER_66_323 ();
 FILLCELL_X1 FILLER_66_352 ();
 FILLCELL_X2 FILLER_66_366 ();
 FILLCELL_X4 FILLER_66_370 ();
 FILLCELL_X2 FILLER_66_374 ();
 FILLCELL_X4 FILLER_66_379 ();
 FILLCELL_X32 FILLER_66_411 ();
 FILLCELL_X4 FILLER_66_443 ();
 FILLCELL_X1 FILLER_66_447 ();
 FILLCELL_X1 FILLER_66_470 ();
 FILLCELL_X2 FILLER_66_487 ();
 FILLCELL_X2 FILLER_66_506 ();
 FILLCELL_X8 FILLER_66_616 ();
 FILLCELL_X4 FILLER_66_624 ();
 FILLCELL_X2 FILLER_66_628 ();
 FILLCELL_X1 FILLER_66_630 ();
 FILLCELL_X2 FILLER_66_646 ();
 FILLCELL_X16 FILLER_66_659 ();
 FILLCELL_X4 FILLER_66_675 ();
 FILLCELL_X1 FILLER_66_720 ();
 FILLCELL_X1 FILLER_66_783 ();
 FILLCELL_X2 FILLER_66_837 ();
 FILLCELL_X1 FILLER_66_849 ();
 FILLCELL_X1 FILLER_66_868 ();
 FILLCELL_X1 FILLER_66_884 ();
 FILLCELL_X2 FILLER_66_925 ();
 FILLCELL_X4 FILLER_66_972 ();
 FILLCELL_X2 FILLER_66_976 ();
 FILLCELL_X2 FILLER_66_1034 ();
 FILLCELL_X1 FILLER_66_1052 ();
 FILLCELL_X4 FILLER_66_1092 ();
 FILLCELL_X4 FILLER_66_1099 ();
 FILLCELL_X8 FILLER_66_1125 ();
 FILLCELL_X1 FILLER_66_1133 ();
 FILLCELL_X4 FILLER_66_1143 ();
 FILLCELL_X1 FILLER_66_1147 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X8 FILLER_67_33 ();
 FILLCELL_X1 FILLER_67_41 ();
 FILLCELL_X1 FILLER_67_71 ();
 FILLCELL_X2 FILLER_67_86 ();
 FILLCELL_X1 FILLER_67_98 ();
 FILLCELL_X1 FILLER_67_103 ();
 FILLCELL_X1 FILLER_67_168 ();
 FILLCELL_X1 FILLER_67_181 ();
 FILLCELL_X1 FILLER_67_186 ();
 FILLCELL_X1 FILLER_67_190 ();
 FILLCELL_X1 FILLER_67_193 ();
 FILLCELL_X4 FILLER_67_209 ();
 FILLCELL_X1 FILLER_67_213 ();
 FILLCELL_X16 FILLER_67_234 ();
 FILLCELL_X1 FILLER_67_250 ();
 FILLCELL_X4 FILLER_67_263 ();
 FILLCELL_X2 FILLER_67_267 ();
 FILLCELL_X1 FILLER_67_269 ();
 FILLCELL_X1 FILLER_67_286 ();
 FILLCELL_X8 FILLER_67_311 ();
 FILLCELL_X2 FILLER_67_319 ();
 FILLCELL_X2 FILLER_67_343 ();
 FILLCELL_X1 FILLER_67_345 ();
 FILLCELL_X2 FILLER_67_353 ();
 FILLCELL_X1 FILLER_67_393 ();
 FILLCELL_X1 FILLER_67_396 ();
 FILLCELL_X1 FILLER_67_399 ();
 FILLCELL_X2 FILLER_67_404 ();
 FILLCELL_X16 FILLER_67_412 ();
 FILLCELL_X4 FILLER_67_428 ();
 FILLCELL_X1 FILLER_67_432 ();
 FILLCELL_X2 FILLER_67_455 ();
 FILLCELL_X2 FILLER_67_499 ();
 FILLCELL_X4 FILLER_67_526 ();
 FILLCELL_X1 FILLER_67_530 ();
 FILLCELL_X1 FILLER_67_558 ();
 FILLCELL_X2 FILLER_67_588 ();
 FILLCELL_X4 FILLER_67_601 ();
 FILLCELL_X1 FILLER_67_605 ();
 FILLCELL_X2 FILLER_67_613 ();
 FILLCELL_X8 FILLER_67_627 ();
 FILLCELL_X4 FILLER_67_635 ();
 FILLCELL_X2 FILLER_67_639 ();
 FILLCELL_X4 FILLER_67_647 ();
 FILLCELL_X1 FILLER_67_651 ();
 FILLCELL_X4 FILLER_67_658 ();
 FILLCELL_X1 FILLER_67_662 ();
 FILLCELL_X16 FILLER_67_666 ();
 FILLCELL_X8 FILLER_67_682 ();
 FILLCELL_X4 FILLER_67_694 ();
 FILLCELL_X1 FILLER_67_728 ();
 FILLCELL_X1 FILLER_67_736 ();
 FILLCELL_X2 FILLER_67_911 ();
 FILLCELL_X1 FILLER_67_1003 ();
 FILLCELL_X2 FILLER_67_1027 ();
 FILLCELL_X1 FILLER_67_1053 ();
 FILLCELL_X16 FILLER_67_1095 ();
 FILLCELL_X4 FILLER_67_1111 ();
 FILLCELL_X1 FILLER_67_1115 ();
 FILLCELL_X2 FILLER_67_1139 ();
 FILLCELL_X1 FILLER_67_1141 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X16 FILLER_68_33 ();
 FILLCELL_X4 FILLER_68_49 ();
 FILLCELL_X1 FILLER_68_53 ();
 FILLCELL_X8 FILLER_68_74 ();
 FILLCELL_X4 FILLER_68_82 ();
 FILLCELL_X2 FILLER_68_86 ();
 FILLCELL_X1 FILLER_68_88 ();
 FILLCELL_X1 FILLER_68_108 ();
 FILLCELL_X2 FILLER_68_111 ();
 FILLCELL_X1 FILLER_68_113 ();
 FILLCELL_X2 FILLER_68_126 ();
 FILLCELL_X1 FILLER_68_128 ();
 FILLCELL_X4 FILLER_68_175 ();
 FILLCELL_X1 FILLER_68_179 ();
 FILLCELL_X2 FILLER_68_213 ();
 FILLCELL_X1 FILLER_68_247 ();
 FILLCELL_X4 FILLER_68_282 ();
 FILLCELL_X1 FILLER_68_295 ();
 FILLCELL_X8 FILLER_68_302 ();
 FILLCELL_X4 FILLER_68_310 ();
 FILLCELL_X4 FILLER_68_324 ();
 FILLCELL_X8 FILLER_68_342 ();
 FILLCELL_X4 FILLER_68_360 ();
 FILLCELL_X2 FILLER_68_373 ();
 FILLCELL_X16 FILLER_68_404 ();
 FILLCELL_X2 FILLER_68_420 ();
 FILLCELL_X1 FILLER_68_422 ();
 FILLCELL_X1 FILLER_68_448 ();
 FILLCELL_X1 FILLER_68_528 ();
 FILLCELL_X1 FILLER_68_556 ();
 FILLCELL_X1 FILLER_68_589 ();
 FILLCELL_X1 FILLER_68_603 ();
 FILLCELL_X1 FILLER_68_619 ();
 FILLCELL_X8 FILLER_68_632 ();
 FILLCELL_X2 FILLER_68_640 ();
 FILLCELL_X1 FILLER_68_642 ();
 FILLCELL_X1 FILLER_68_646 ();
 FILLCELL_X16 FILLER_68_653 ();
 FILLCELL_X4 FILLER_68_669 ();
 FILLCELL_X2 FILLER_68_673 ();
 FILLCELL_X1 FILLER_68_695 ();
 FILLCELL_X1 FILLER_68_798 ();
 FILLCELL_X1 FILLER_68_859 ();
 FILLCELL_X2 FILLER_68_936 ();
 FILLCELL_X1 FILLER_68_938 ();
 FILLCELL_X1 FILLER_68_963 ();
 FILLCELL_X1 FILLER_68_971 ();
 FILLCELL_X1 FILLER_68_976 ();
 FILLCELL_X4 FILLER_68_998 ();
 FILLCELL_X1 FILLER_68_1020 ();
 FILLCELL_X1 FILLER_68_1025 ();
 FILLCELL_X2 FILLER_68_1035 ();
 FILLCELL_X1 FILLER_68_1052 ();
 FILLCELL_X1 FILLER_68_1055 ();
 FILLCELL_X1 FILLER_68_1066 ();
 FILLCELL_X8 FILLER_68_1080 ();
 FILLCELL_X1 FILLER_68_1099 ();
 FILLCELL_X1 FILLER_68_1103 ();
 FILLCELL_X1 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X8 FILLER_69_33 ();
 FILLCELL_X4 FILLER_69_41 ();
 FILLCELL_X1 FILLER_69_45 ();
 FILLCELL_X1 FILLER_69_96 ();
 FILLCELL_X2 FILLER_69_103 ();
 FILLCELL_X1 FILLER_69_107 ();
 FILLCELL_X4 FILLER_69_145 ();
 FILLCELL_X2 FILLER_69_149 ();
 FILLCELL_X2 FILLER_69_153 ();
 FILLCELL_X1 FILLER_69_199 ();
 FILLCELL_X8 FILLER_69_206 ();
 FILLCELL_X4 FILLER_69_261 ();
 FILLCELL_X1 FILLER_69_268 ();
 FILLCELL_X1 FILLER_69_286 ();
 FILLCELL_X2 FILLER_69_291 ();
 FILLCELL_X1 FILLER_69_293 ();
 FILLCELL_X2 FILLER_69_319 ();
 FILLCELL_X8 FILLER_69_335 ();
 FILLCELL_X2 FILLER_69_409 ();
 FILLCELL_X1 FILLER_69_413 ();
 FILLCELL_X1 FILLER_69_434 ();
 FILLCELL_X1 FILLER_69_442 ();
 FILLCELL_X1 FILLER_69_450 ();
 FILLCELL_X1 FILLER_69_476 ();
 FILLCELL_X1 FILLER_69_480 ();
 FILLCELL_X2 FILLER_69_498 ();
 FILLCELL_X1 FILLER_69_580 ();
 FILLCELL_X1 FILLER_69_585 ();
 FILLCELL_X8 FILLER_69_624 ();
 FILLCELL_X32 FILLER_69_639 ();
 FILLCELL_X2 FILLER_69_671 ();
 FILLCELL_X1 FILLER_69_689 ();
 FILLCELL_X1 FILLER_69_697 ();
 FILLCELL_X1 FILLER_69_706 ();
 FILLCELL_X1 FILLER_69_728 ();
 FILLCELL_X2 FILLER_69_996 ();
 FILLCELL_X1 FILLER_69_998 ();
 FILLCELL_X2 FILLER_69_1005 ();
 FILLCELL_X1 FILLER_69_1007 ();
 FILLCELL_X1 FILLER_69_1012 ();
 FILLCELL_X2 FILLER_69_1016 ();
 FILLCELL_X1 FILLER_69_1018 ();
 FILLCELL_X2 FILLER_69_1023 ();
 FILLCELL_X1 FILLER_69_1025 ();
 FILLCELL_X2 FILLER_69_1035 ();
 FILLCELL_X1 FILLER_69_1037 ();
 FILLCELL_X4 FILLER_69_1079 ();
 FILLCELL_X1 FILLER_69_1090 ();
 FILLCELL_X2 FILLER_69_1146 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X2 FILLER_70_103 ();
 FILLCELL_X1 FILLER_70_105 ();
 FILLCELL_X16 FILLER_70_113 ();
 FILLCELL_X8 FILLER_70_129 ();
 FILLCELL_X2 FILLER_70_137 ();
 FILLCELL_X1 FILLER_70_139 ();
 FILLCELL_X2 FILLER_70_153 ();
 FILLCELL_X1 FILLER_70_155 ();
 FILLCELL_X4 FILLER_70_191 ();
 FILLCELL_X4 FILLER_70_216 ();
 FILLCELL_X2 FILLER_70_220 ();
 FILLCELL_X1 FILLER_70_222 ();
 FILLCELL_X2 FILLER_70_226 ();
 FILLCELL_X1 FILLER_70_228 ();
 FILLCELL_X2 FILLER_70_246 ();
 FILLCELL_X2 FILLER_70_270 ();
 FILLCELL_X2 FILLER_70_278 ();
 FILLCELL_X1 FILLER_70_280 ();
 FILLCELL_X2 FILLER_70_285 ();
 FILLCELL_X2 FILLER_70_301 ();
 FILLCELL_X1 FILLER_70_308 ();
 FILLCELL_X1 FILLER_70_318 ();
 FILLCELL_X2 FILLER_70_321 ();
 FILLCELL_X1 FILLER_70_329 ();
 FILLCELL_X1 FILLER_70_349 ();
 FILLCELL_X2 FILLER_70_362 ();
 FILLCELL_X1 FILLER_70_364 ();
 FILLCELL_X2 FILLER_70_368 ();
 FILLCELL_X2 FILLER_70_382 ();
 FILLCELL_X1 FILLER_70_384 ();
 FILLCELL_X8 FILLER_70_389 ();
 FILLCELL_X4 FILLER_70_397 ();
 FILLCELL_X2 FILLER_70_401 ();
 FILLCELL_X1 FILLER_70_403 ();
 FILLCELL_X4 FILLER_70_416 ();
 FILLCELL_X2 FILLER_70_420 ();
 FILLCELL_X1 FILLER_70_434 ();
 FILLCELL_X4 FILLER_70_442 ();
 FILLCELL_X1 FILLER_70_488 ();
 FILLCELL_X2 FILLER_70_534 ();
 FILLCELL_X1 FILLER_70_594 ();
 FILLCELL_X1 FILLER_70_598 ();
 FILLCELL_X1 FILLER_70_603 ();
 FILLCELL_X2 FILLER_70_620 ();
 FILLCELL_X1 FILLER_70_622 ();
 FILLCELL_X2 FILLER_70_628 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X16 FILLER_70_637 ();
 FILLCELL_X8 FILLER_70_653 ();
 FILLCELL_X1 FILLER_70_661 ();
 FILLCELL_X1 FILLER_70_684 ();
 FILLCELL_X1 FILLER_70_692 ();
 FILLCELL_X1 FILLER_70_700 ();
 FILLCELL_X1 FILLER_70_706 ();
 FILLCELL_X2 FILLER_70_773 ();
 FILLCELL_X1 FILLER_70_880 ();
 FILLCELL_X2 FILLER_70_939 ();
 FILLCELL_X2 FILLER_70_969 ();
 FILLCELL_X1 FILLER_70_982 ();
 FILLCELL_X1 FILLER_70_986 ();
 FILLCELL_X1 FILLER_70_992 ();
 FILLCELL_X1 FILLER_70_997 ();
 FILLCELL_X2 FILLER_70_1018 ();
 FILLCELL_X4 FILLER_70_1033 ();
 FILLCELL_X2 FILLER_70_1037 ();
 FILLCELL_X1 FILLER_70_1039 ();
 FILLCELL_X4 FILLER_70_1044 ();
 FILLCELL_X2 FILLER_70_1048 ();
 FILLCELL_X1 FILLER_70_1058 ();
 FILLCELL_X1 FILLER_70_1062 ();
 FILLCELL_X2 FILLER_70_1071 ();
 FILLCELL_X2 FILLER_70_1126 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X4 FILLER_71_33 ();
 FILLCELL_X16 FILLER_71_43 ();
 FILLCELL_X2 FILLER_71_59 ();
 FILLCELL_X1 FILLER_71_61 ();
 FILLCELL_X8 FILLER_71_65 ();
 FILLCELL_X4 FILLER_71_73 ();
 FILLCELL_X1 FILLER_71_77 ();
 FILLCELL_X1 FILLER_71_100 ();
 FILLCELL_X4 FILLER_71_117 ();
 FILLCELL_X4 FILLER_71_123 ();
 FILLCELL_X2 FILLER_71_169 ();
 FILLCELL_X2 FILLER_71_185 ();
 FILLCELL_X1 FILLER_71_191 ();
 FILLCELL_X1 FILLER_71_202 ();
 FILLCELL_X4 FILLER_71_208 ();
 FILLCELL_X2 FILLER_71_212 ();
 FILLCELL_X1 FILLER_71_247 ();
 FILLCELL_X2 FILLER_71_255 ();
 FILLCELL_X1 FILLER_71_276 ();
 FILLCELL_X1 FILLER_71_280 ();
 FILLCELL_X1 FILLER_71_301 ();
 FILLCELL_X2 FILLER_71_322 ();
 FILLCELL_X2 FILLER_71_341 ();
 FILLCELL_X1 FILLER_71_343 ();
 FILLCELL_X32 FILLER_71_354 ();
 FILLCELL_X4 FILLER_71_386 ();
 FILLCELL_X2 FILLER_71_390 ();
 FILLCELL_X1 FILLER_71_392 ();
 FILLCELL_X8 FILLER_71_423 ();
 FILLCELL_X1 FILLER_71_445 ();
 FILLCELL_X1 FILLER_71_608 ();
 FILLCELL_X16 FILLER_71_656 ();
 FILLCELL_X4 FILLER_71_672 ();
 FILLCELL_X2 FILLER_71_676 ();
 FILLCELL_X2 FILLER_71_698 ();
 FILLCELL_X1 FILLER_71_727 ();
 FILLCELL_X1 FILLER_71_736 ();
 FILLCELL_X1 FILLER_71_780 ();
 FILLCELL_X1 FILLER_71_836 ();
 FILLCELL_X1 FILLER_71_898 ();
 FILLCELL_X2 FILLER_71_987 ();
 FILLCELL_X2 FILLER_71_1029 ();
 FILLCELL_X2 FILLER_71_1042 ();
 FILLCELL_X2 FILLER_71_1061 ();
 FILLCELL_X1 FILLER_71_1071 ();
 FILLCELL_X1 FILLER_71_1082 ();
 FILLCELL_X1 FILLER_71_1122 ();
 FILLCELL_X1 FILLER_72_1 ();
 FILLCELL_X4 FILLER_72_25 ();
 FILLCELL_X4 FILLER_72_31 ();
 FILLCELL_X2 FILLER_72_35 ();
 FILLCELL_X4 FILLER_72_89 ();
 FILLCELL_X2 FILLER_72_93 ();
 FILLCELL_X2 FILLER_72_97 ();
 FILLCELL_X1 FILLER_72_99 ();
 FILLCELL_X8 FILLER_72_124 ();
 FILLCELL_X4 FILLER_72_152 ();
 FILLCELL_X2 FILLER_72_156 ();
 FILLCELL_X1 FILLER_72_158 ();
 FILLCELL_X1 FILLER_72_172 ();
 FILLCELL_X1 FILLER_72_193 ();
 FILLCELL_X1 FILLER_72_224 ();
 FILLCELL_X2 FILLER_72_256 ();
 FILLCELL_X1 FILLER_72_289 ();
 FILLCELL_X2 FILLER_72_333 ();
 FILLCELL_X4 FILLER_72_337 ();
 FILLCELL_X32 FILLER_72_351 ();
 FILLCELL_X8 FILLER_72_383 ();
 FILLCELL_X2 FILLER_72_391 ();
 FILLCELL_X1 FILLER_72_393 ();
 FILLCELL_X2 FILLER_72_416 ();
 FILLCELL_X2 FILLER_72_425 ();
 FILLCELL_X4 FILLER_72_434 ();
 FILLCELL_X1 FILLER_72_545 ();
 FILLCELL_X1 FILLER_72_573 ();
 FILLCELL_X1 FILLER_72_587 ();
 FILLCELL_X1 FILLER_72_592 ();
 FILLCELL_X1 FILLER_72_596 ();
 FILLCELL_X2 FILLER_72_613 ();
 FILLCELL_X8 FILLER_72_652 ();
 FILLCELL_X2 FILLER_72_680 ();
 FILLCELL_X1 FILLER_72_684 ();
 FILLCELL_X4 FILLER_72_687 ();
 FILLCELL_X1 FILLER_72_698 ();
 FILLCELL_X1 FILLER_72_706 ();
 FILLCELL_X1 FILLER_72_740 ();
 FILLCELL_X2 FILLER_72_767 ();
 FILLCELL_X1 FILLER_72_796 ();
 FILLCELL_X1 FILLER_72_916 ();
 FILLCELL_X1 FILLER_72_957 ();
 FILLCELL_X1 FILLER_72_963 ();
 FILLCELL_X1 FILLER_72_972 ();
 FILLCELL_X1 FILLER_72_980 ();
 FILLCELL_X1 FILLER_72_1001 ();
 FILLCELL_X1 FILLER_72_1016 ();
 FILLCELL_X1 FILLER_72_1046 ();
 FILLCELL_X1 FILLER_72_1051 ();
 FILLCELL_X1 FILLER_72_1055 ();
 FILLCELL_X2 FILLER_72_1060 ();
 FILLCELL_X1 FILLER_72_1093 ();
 FILLCELL_X1 FILLER_72_1101 ();
 FILLCELL_X2 FILLER_72_1121 ();
 FILLCELL_X1 FILLER_72_1127 ();
 FILLCELL_X2 FILLER_73_5 ();
 FILLCELL_X2 FILLER_73_41 ();
 FILLCELL_X1 FILLER_73_47 ();
 FILLCELL_X4 FILLER_73_67 ();
 FILLCELL_X2 FILLER_73_71 ();
 FILLCELL_X1 FILLER_73_73 ();
 FILLCELL_X1 FILLER_73_85 ();
 FILLCELL_X1 FILLER_73_118 ();
 FILLCELL_X4 FILLER_73_146 ();
 FILLCELL_X1 FILLER_73_210 ();
 FILLCELL_X1 FILLER_73_215 ();
 FILLCELL_X1 FILLER_73_220 ();
 FILLCELL_X4 FILLER_73_250 ();
 FILLCELL_X2 FILLER_73_254 ();
 FILLCELL_X1 FILLER_73_256 ();
 FILLCELL_X2 FILLER_73_259 ();
 FILLCELL_X1 FILLER_73_261 ();
 FILLCELL_X4 FILLER_73_267 ();
 FILLCELL_X8 FILLER_73_281 ();
 FILLCELL_X2 FILLER_73_289 ();
 FILLCELL_X1 FILLER_73_291 ();
 FILLCELL_X8 FILLER_73_305 ();
 FILLCELL_X2 FILLER_73_313 ();
 FILLCELL_X1 FILLER_73_315 ();
 FILLCELL_X2 FILLER_73_352 ();
 FILLCELL_X32 FILLER_73_360 ();
 FILLCELL_X1 FILLER_73_392 ();
 FILLCELL_X4 FILLER_73_415 ();
 FILLCELL_X2 FILLER_73_426 ();
 FILLCELL_X4 FILLER_73_437 ();
 FILLCELL_X2 FILLER_73_441 ();
 FILLCELL_X1 FILLER_73_466 ();
 FILLCELL_X2 FILLER_73_495 ();
 FILLCELL_X1 FILLER_73_531 ();
 FILLCELL_X2 FILLER_73_563 ();
 FILLCELL_X1 FILLER_73_574 ();
 FILLCELL_X1 FILLER_73_582 ();
 FILLCELL_X1 FILLER_73_586 ();
 FILLCELL_X1 FILLER_73_633 ();
 FILLCELL_X1 FILLER_73_653 ();
 FILLCELL_X8 FILLER_73_663 ();
 FILLCELL_X2 FILLER_73_714 ();
 FILLCELL_X1 FILLER_73_775 ();
 FILLCELL_X1 FILLER_73_779 ();
 FILLCELL_X1 FILLER_73_935 ();
 FILLCELL_X1 FILLER_73_960 ();
 FILLCELL_X2 FILLER_73_982 ();
 FILLCELL_X1 FILLER_73_1008 ();
 FILLCELL_X1 FILLER_73_1016 ();
 FILLCELL_X1 FILLER_73_1023 ();
 FILLCELL_X1 FILLER_73_1034 ();
 FILLCELL_X2 FILLER_73_1040 ();
 FILLCELL_X2 FILLER_73_1046 ();
 FILLCELL_X1 FILLER_73_1052 ();
 FILLCELL_X2 FILLER_73_1060 ();
 FILLCELL_X2 FILLER_73_1124 ();
 FILLCELL_X4 FILLER_74_20 ();
 FILLCELL_X2 FILLER_74_24 ();
 FILLCELL_X1 FILLER_74_26 ();
 FILLCELL_X2 FILLER_74_61 ();
 FILLCELL_X1 FILLER_74_63 ();
 FILLCELL_X8 FILLER_74_66 ();
 FILLCELL_X4 FILLER_74_74 ();
 FILLCELL_X8 FILLER_74_142 ();
 FILLCELL_X2 FILLER_74_150 ();
 FILLCELL_X2 FILLER_74_156 ();
 FILLCELL_X1 FILLER_74_158 ();
 FILLCELL_X1 FILLER_74_163 ();
 FILLCELL_X4 FILLER_74_175 ();
 FILLCELL_X1 FILLER_74_181 ();
 FILLCELL_X2 FILLER_74_212 ();
 FILLCELL_X1 FILLER_74_228 ();
 FILLCELL_X1 FILLER_74_247 ();
 FILLCELL_X1 FILLER_74_252 ();
 FILLCELL_X8 FILLER_74_263 ();
 FILLCELL_X1 FILLER_74_271 ();
 FILLCELL_X2 FILLER_74_277 ();
 FILLCELL_X1 FILLER_74_279 ();
 FILLCELL_X2 FILLER_74_294 ();
 FILLCELL_X2 FILLER_74_300 ();
 FILLCELL_X1 FILLER_74_302 ();
 FILLCELL_X1 FILLER_74_321 ();
 FILLCELL_X2 FILLER_74_332 ();
 FILLCELL_X2 FILLER_74_346 ();
 FILLCELL_X1 FILLER_74_348 ();
 FILLCELL_X16 FILLER_74_353 ();
 FILLCELL_X2 FILLER_74_369 ();
 FILLCELL_X16 FILLER_74_379 ();
 FILLCELL_X2 FILLER_74_395 ();
 FILLCELL_X1 FILLER_74_463 ();
 FILLCELL_X1 FILLER_74_577 ();
 FILLCELL_X1 FILLER_74_587 ();
 FILLCELL_X2 FILLER_74_619 ();
 FILLCELL_X1 FILLER_74_621 ();
 FILLCELL_X32 FILLER_74_658 ();
 FILLCELL_X1 FILLER_74_898 ();
 FILLCELL_X1 FILLER_74_902 ();
 FILLCELL_X1 FILLER_74_923 ();
 FILLCELL_X1 FILLER_74_934 ();
 FILLCELL_X1 FILLER_74_955 ();
 FILLCELL_X1 FILLER_74_960 ();
 FILLCELL_X1 FILLER_74_968 ();
 FILLCELL_X1 FILLER_74_973 ();
 FILLCELL_X8 FILLER_74_978 ();
 FILLCELL_X4 FILLER_74_986 ();
 FILLCELL_X1 FILLER_74_999 ();
 FILLCELL_X1 FILLER_74_1029 ();
 FILLCELL_X1 FILLER_74_1057 ();
 FILLCELL_X4 FILLER_74_1138 ();
 FILLCELL_X4 FILLER_75_4 ();
 FILLCELL_X1 FILLER_75_11 ();
 FILLCELL_X1 FILLER_75_53 ();
 FILLCELL_X4 FILLER_75_112 ();
 FILLCELL_X1 FILLER_75_140 ();
 FILLCELL_X2 FILLER_75_153 ();
 FILLCELL_X2 FILLER_75_157 ();
 FILLCELL_X4 FILLER_75_207 ();
 FILLCELL_X1 FILLER_75_211 ();
 FILLCELL_X1 FILLER_75_266 ();
 FILLCELL_X2 FILLER_75_270 ();
 FILLCELL_X1 FILLER_75_282 ();
 FILLCELL_X4 FILLER_75_293 ();
 FILLCELL_X1 FILLER_75_297 ();
 FILLCELL_X8 FILLER_75_304 ();
 FILLCELL_X4 FILLER_75_312 ();
 FILLCELL_X1 FILLER_75_316 ();
 FILLCELL_X1 FILLER_75_327 ();
 FILLCELL_X2 FILLER_75_348 ();
 FILLCELL_X32 FILLER_75_354 ();
 FILLCELL_X4 FILLER_75_386 ();
 FILLCELL_X2 FILLER_75_390 ();
 FILLCELL_X1 FILLER_75_392 ();
 FILLCELL_X2 FILLER_75_415 ();
 FILLCELL_X2 FILLER_75_446 ();
 FILLCELL_X2 FILLER_75_451 ();
 FILLCELL_X1 FILLER_75_654 ();
 FILLCELL_X16 FILLER_75_658 ();
 FILLCELL_X2 FILLER_75_674 ();
 FILLCELL_X1 FILLER_75_696 ();
 FILLCELL_X2 FILLER_75_746 ();
 FILLCELL_X1 FILLER_75_748 ();
 FILLCELL_X1 FILLER_75_784 ();
 FILLCELL_X1 FILLER_75_970 ();
 FILLCELL_X16 FILLER_75_978 ();
 FILLCELL_X1 FILLER_75_994 ();
 FILLCELL_X8 FILLER_75_1035 ();
 FILLCELL_X1 FILLER_75_1043 ();
 FILLCELL_X4 FILLER_75_1053 ();
 FILLCELL_X1 FILLER_75_1125 ();
 FILLCELL_X8 FILLER_76_7 ();
 FILLCELL_X4 FILLER_76_15 ();
 FILLCELL_X1 FILLER_76_19 ();
 FILLCELL_X4 FILLER_76_22 ();
 FILLCELL_X8 FILLER_76_60 ();
 FILLCELL_X2 FILLER_76_68 ();
 FILLCELL_X1 FILLER_76_70 ();
 FILLCELL_X2 FILLER_76_75 ();
 FILLCELL_X1 FILLER_76_77 ();
 FILLCELL_X4 FILLER_76_148 ();
 FILLCELL_X8 FILLER_76_172 ();
 FILLCELL_X4 FILLER_76_180 ();
 FILLCELL_X4 FILLER_76_194 ();
 FILLCELL_X2 FILLER_76_198 ();
 FILLCELL_X2 FILLER_76_249 ();
 FILLCELL_X1 FILLER_76_267 ();
 FILLCELL_X4 FILLER_76_279 ();
 FILLCELL_X16 FILLER_76_294 ();
 FILLCELL_X8 FILLER_76_310 ();
 FILLCELL_X4 FILLER_76_318 ();
 FILLCELL_X1 FILLER_76_322 ();
 FILLCELL_X2 FILLER_76_329 ();
 FILLCELL_X4 FILLER_76_337 ();
 FILLCELL_X2 FILLER_76_341 ();
 FILLCELL_X32 FILLER_76_345 ();
 FILLCELL_X8 FILLER_76_377 ();
 FILLCELL_X4 FILLER_76_385 ();
 FILLCELL_X1 FILLER_76_389 ();
 FILLCELL_X2 FILLER_76_410 ();
 FILLCELL_X1 FILLER_76_436 ();
 FILLCELL_X1 FILLER_76_443 ();
 FILLCELL_X2 FILLER_76_532 ();
 FILLCELL_X1 FILLER_76_588 ();
 FILLCELL_X1 FILLER_76_602 ();
 FILLCELL_X1 FILLER_76_630 ();
 FILLCELL_X2 FILLER_76_645 ();
 FILLCELL_X32 FILLER_76_652 ();
 FILLCELL_X8 FILLER_76_684 ();
 FILLCELL_X1 FILLER_76_692 ();
 FILLCELL_X2 FILLER_76_767 ();
 FILLCELL_X2 FILLER_76_854 ();
 FILLCELL_X1 FILLER_76_872 ();
 FILLCELL_X1 FILLER_76_920 ();
 FILLCELL_X1 FILLER_76_945 ();
 FILLCELL_X4 FILLER_76_969 ();
 FILLCELL_X1 FILLER_76_973 ();
 FILLCELL_X2 FILLER_76_995 ();
 FILLCELL_X1 FILLER_76_1009 ();
 FILLCELL_X2 FILLER_76_1041 ();
 FILLCELL_X1 FILLER_76_1043 ();
 FILLCELL_X2 FILLER_76_1116 ();
 FILLCELL_X1 FILLER_76_1118 ();
 FILLCELL_X2 FILLER_76_1143 ();
 FILLCELL_X1 FILLER_77_13 ();
 FILLCELL_X2 FILLER_77_50 ();
 FILLCELL_X4 FILLER_77_84 ();
 FILLCELL_X2 FILLER_77_88 ();
 FILLCELL_X4 FILLER_77_92 ();
 FILLCELL_X8 FILLER_77_138 ();
 FILLCELL_X1 FILLER_77_146 ();
 FILLCELL_X1 FILLER_77_153 ();
 FILLCELL_X2 FILLER_77_162 ();
 FILLCELL_X16 FILLER_77_186 ();
 FILLCELL_X8 FILLER_77_202 ();
 FILLCELL_X4 FILLER_77_210 ();
 FILLCELL_X2 FILLER_77_214 ();
 FILLCELL_X1 FILLER_77_237 ();
 FILLCELL_X1 FILLER_77_242 ();
 FILLCELL_X4 FILLER_77_264 ();
 FILLCELL_X4 FILLER_77_290 ();
 FILLCELL_X2 FILLER_77_294 ();
 FILLCELL_X2 FILLER_77_326 ();
 FILLCELL_X2 FILLER_77_338 ();
 FILLCELL_X1 FILLER_77_340 ();
 FILLCELL_X1 FILLER_77_357 ();
 FILLCELL_X16 FILLER_77_368 ();
 FILLCELL_X4 FILLER_77_384 ();
 FILLCELL_X2 FILLER_77_410 ();
 FILLCELL_X1 FILLER_77_412 ();
 FILLCELL_X1 FILLER_77_423 ();
 FILLCELL_X1 FILLER_77_565 ();
 FILLCELL_X1 FILLER_77_587 ();
 FILLCELL_X2 FILLER_77_629 ();
 FILLCELL_X4 FILLER_77_646 ();
 FILLCELL_X2 FILLER_77_650 ();
 FILLCELL_X16 FILLER_77_657 ();
 FILLCELL_X4 FILLER_77_673 ();
 FILLCELL_X1 FILLER_77_728 ();
 FILLCELL_X1 FILLER_77_880 ();
 FILLCELL_X2 FILLER_77_885 ();
 FILLCELL_X1 FILLER_77_907 ();
 FILLCELL_X2 FILLER_77_914 ();
 FILLCELL_X1 FILLER_77_920 ();
 FILLCELL_X2 FILLER_77_925 ();
 FILLCELL_X4 FILLER_77_949 ();
 FILLCELL_X1 FILLER_77_953 ();
 FILLCELL_X2 FILLER_77_964 ();
 FILLCELL_X1 FILLER_77_996 ();
 FILLCELL_X4 FILLER_77_1013 ();
 FILLCELL_X1 FILLER_77_1040 ();
 FILLCELL_X1 FILLER_77_1045 ();
 FILLCELL_X1 FILLER_77_1066 ();
 FILLCELL_X2 FILLER_78_31 ();
 FILLCELL_X4 FILLER_78_37 ();
 FILLCELL_X1 FILLER_78_41 ();
 FILLCELL_X2 FILLER_78_44 ();
 FILLCELL_X1 FILLER_78_46 ();
 FILLCELL_X2 FILLER_78_53 ();
 FILLCELL_X1 FILLER_78_55 ();
 FILLCELL_X4 FILLER_78_140 ();
 FILLCELL_X2 FILLER_78_144 ();
 FILLCELL_X1 FILLER_78_146 ();
 FILLCELL_X1 FILLER_78_157 ();
 FILLCELL_X1 FILLER_78_169 ();
 FILLCELL_X8 FILLER_78_209 ();
 FILLCELL_X2 FILLER_78_217 ();
 FILLCELL_X1 FILLER_78_223 ();
 FILLCELL_X2 FILLER_78_232 ();
 FILLCELL_X1 FILLER_78_234 ();
 FILLCELL_X4 FILLER_78_245 ();
 FILLCELL_X4 FILLER_78_263 ();
 FILLCELL_X16 FILLER_78_307 ();
 FILLCELL_X1 FILLER_78_346 ();
 FILLCELL_X2 FILLER_78_353 ();
 FILLCELL_X1 FILLER_78_355 ();
 FILLCELL_X32 FILLER_78_362 ();
 FILLCELL_X4 FILLER_78_394 ();
 FILLCELL_X2 FILLER_78_398 ();
 FILLCELL_X1 FILLER_78_400 ();
 FILLCELL_X2 FILLER_78_426 ();
 FILLCELL_X4 FILLER_78_431 ();
 FILLCELL_X2 FILLER_78_441 ();
 FILLCELL_X1 FILLER_78_522 ();
 FILLCELL_X1 FILLER_78_574 ();
 FILLCELL_X1 FILLER_78_614 ();
 FILLCELL_X32 FILLER_78_650 ();
 FILLCELL_X8 FILLER_78_682 ();
 FILLCELL_X2 FILLER_78_692 ();
 FILLCELL_X1 FILLER_78_869 ();
 FILLCELL_X1 FILLER_78_902 ();
 FILLCELL_X2 FILLER_78_954 ();
 FILLCELL_X1 FILLER_78_956 ();
 FILLCELL_X1 FILLER_78_975 ();
 FILLCELL_X2 FILLER_78_990 ();
 FILLCELL_X1 FILLER_78_1018 ();
 FILLCELL_X2 FILLER_78_1029 ();
 FILLCELL_X1 FILLER_78_1071 ();
 FILLCELL_X1 FILLER_78_1077 ();
 FILLCELL_X1 FILLER_78_1081 ();
 FILLCELL_X1 FILLER_78_1132 ();
 FILLCELL_X2 FILLER_78_1145 ();
 FILLCELL_X1 FILLER_78_1147 ();
 FILLCELL_X8 FILLER_79_58 ();
 FILLCELL_X1 FILLER_79_87 ();
 FILLCELL_X8 FILLER_79_104 ();
 FILLCELL_X1 FILLER_79_112 ();
 FILLCELL_X16 FILLER_79_115 ();
 FILLCELL_X4 FILLER_79_131 ();
 FILLCELL_X2 FILLER_79_135 ();
 FILLCELL_X8 FILLER_79_139 ();
 FILLCELL_X4 FILLER_79_147 ();
 FILLCELL_X2 FILLER_79_151 ();
 FILLCELL_X4 FILLER_79_200 ();
 FILLCELL_X4 FILLER_79_214 ();
 FILLCELL_X1 FILLER_79_220 ();
 FILLCELL_X2 FILLER_79_260 ();
 FILLCELL_X2 FILLER_79_284 ();
 FILLCELL_X2 FILLER_79_289 ();
 FILLCELL_X1 FILLER_79_328 ();
 FILLCELL_X2 FILLER_79_345 ();
 FILLCELL_X1 FILLER_79_349 ();
 FILLCELL_X32 FILLER_79_368 ();
 FILLCELL_X16 FILLER_79_400 ();
 FILLCELL_X1 FILLER_79_642 ();
 FILLCELL_X32 FILLER_79_648 ();
 FILLCELL_X16 FILLER_79_680 ();
 FILLCELL_X2 FILLER_79_709 ();
 FILLCELL_X1 FILLER_79_711 ();
 FILLCELL_X2 FILLER_79_714 ();
 FILLCELL_X8 FILLER_79_737 ();
 FILLCELL_X4 FILLER_79_745 ();
 FILLCELL_X1 FILLER_79_749 ();
 FILLCELL_X2 FILLER_79_832 ();
 FILLCELL_X1 FILLER_79_834 ();
 FILLCELL_X2 FILLER_79_868 ();
 FILLCELL_X1 FILLER_79_870 ();
 FILLCELL_X4 FILLER_79_897 ();
 FILLCELL_X2 FILLER_79_905 ();
 FILLCELL_X1 FILLER_79_907 ();
 FILLCELL_X2 FILLER_79_915 ();
 FILLCELL_X1 FILLER_79_917 ();
 FILLCELL_X8 FILLER_79_938 ();
 FILLCELL_X1 FILLER_79_946 ();
 FILLCELL_X8 FILLER_79_994 ();
 FILLCELL_X2 FILLER_79_1002 ();
 FILLCELL_X2 FILLER_79_1146 ();
 FILLCELL_X2 FILLER_80_10 ();
 FILLCELL_X1 FILLER_80_12 ();
 FILLCELL_X1 FILLER_80_20 ();
 FILLCELL_X4 FILLER_80_40 ();
 FILLCELL_X4 FILLER_80_52 ();
 FILLCELL_X2 FILLER_80_56 ();
 FILLCELL_X1 FILLER_80_81 ();
 FILLCELL_X1 FILLER_80_86 ();
 FILLCELL_X1 FILLER_80_94 ();
 FILLCELL_X2 FILLER_80_185 ();
 FILLCELL_X4 FILLER_80_189 ();
 FILLCELL_X2 FILLER_80_193 ();
 FILLCELL_X1 FILLER_80_195 ();
 FILLCELL_X2 FILLER_80_206 ();
 FILLCELL_X8 FILLER_80_212 ();
 FILLCELL_X8 FILLER_80_262 ();
 FILLCELL_X1 FILLER_80_270 ();
 FILLCELL_X4 FILLER_80_293 ();
 FILLCELL_X2 FILLER_80_297 ();
 FILLCELL_X4 FILLER_80_341 ();
 FILLCELL_X4 FILLER_80_357 ();
 FILLCELL_X1 FILLER_80_361 ();
 FILLCELL_X16 FILLER_80_370 ();
 FILLCELL_X1 FILLER_80_386 ();
 FILLCELL_X1 FILLER_80_507 ();
 FILLCELL_X2 FILLER_80_537 ();
 FILLCELL_X1 FILLER_80_571 ();
 FILLCELL_X1 FILLER_80_577 ();
 FILLCELL_X8 FILLER_80_583 ();
 FILLCELL_X4 FILLER_80_591 ();
 FILLCELL_X1 FILLER_80_613 ();
 FILLCELL_X32 FILLER_80_648 ();
 FILLCELL_X16 FILLER_80_680 ();
 FILLCELL_X8 FILLER_80_696 ();
 FILLCELL_X2 FILLER_80_704 ();
 FILLCELL_X4 FILLER_80_722 ();
 FILLCELL_X1 FILLER_80_761 ();
 FILLCELL_X1 FILLER_80_825 ();
 FILLCELL_X4 FILLER_80_835 ();
 FILLCELL_X2 FILLER_80_839 ();
 FILLCELL_X2 FILLER_80_843 ();
 FILLCELL_X1 FILLER_80_845 ();
 FILLCELL_X2 FILLER_80_862 ();
 FILLCELL_X2 FILLER_80_886 ();
 FILLCELL_X1 FILLER_80_919 ();
 FILLCELL_X1 FILLER_80_949 ();
 FILLCELL_X1 FILLER_80_952 ();
 FILLCELL_X1 FILLER_80_957 ();
 FILLCELL_X1 FILLER_80_962 ();
 FILLCELL_X2 FILLER_80_967 ();
 FILLCELL_X1 FILLER_80_969 ();
 FILLCELL_X2 FILLER_80_1015 ();
 FILLCELL_X1 FILLER_80_1017 ();
 FILLCELL_X2 FILLER_80_1047 ();
 FILLCELL_X2 FILLER_80_1063 ();
 FILLCELL_X8 FILLER_81_41 ();
 FILLCELL_X2 FILLER_81_67 ();
 FILLCELL_X1 FILLER_81_69 ();
 FILLCELL_X4 FILLER_81_97 ();
 FILLCELL_X1 FILLER_81_101 ();
 FILLCELL_X1 FILLER_81_122 ();
 FILLCELL_X4 FILLER_81_139 ();
 FILLCELL_X2 FILLER_81_143 ();
 FILLCELL_X1 FILLER_81_168 ();
 FILLCELL_X4 FILLER_81_219 ();
 FILLCELL_X1 FILLER_81_230 ();
 FILLCELL_X1 FILLER_81_240 ();
 FILLCELL_X1 FILLER_81_293 ();
 FILLCELL_X1 FILLER_81_314 ();
 FILLCELL_X1 FILLER_81_348 ();
 FILLCELL_X4 FILLER_81_353 ();
 FILLCELL_X2 FILLER_81_357 ();
 FILLCELL_X1 FILLER_81_365 ();
 FILLCELL_X8 FILLER_81_400 ();
 FILLCELL_X1 FILLER_81_408 ();
 FILLCELL_X1 FILLER_81_413 ();
 FILLCELL_X2 FILLER_81_479 ();
 FILLCELL_X1 FILLER_81_485 ();
 FILLCELL_X2 FILLER_81_491 ();
 FILLCELL_X1 FILLER_81_493 ();
 FILLCELL_X2 FILLER_81_504 ();
 FILLCELL_X1 FILLER_81_506 ();
 FILLCELL_X2 FILLER_81_534 ();
 FILLCELL_X1 FILLER_81_557 ();
 FILLCELL_X1 FILLER_81_564 ();
 FILLCELL_X1 FILLER_81_571 ();
 FILLCELL_X2 FILLER_81_613 ();
 FILLCELL_X2 FILLER_81_632 ();
 FILLCELL_X1 FILLER_81_634 ();
 FILLCELL_X16 FILLER_81_648 ();
 FILLCELL_X8 FILLER_81_664 ();
 FILLCELL_X1 FILLER_81_686 ();
 FILLCELL_X8 FILLER_81_689 ();
 FILLCELL_X4 FILLER_81_697 ();
 FILLCELL_X2 FILLER_81_701 ();
 FILLCELL_X1 FILLER_81_703 ();
 FILLCELL_X1 FILLER_81_748 ();
 FILLCELL_X1 FILLER_81_758 ();
 FILLCELL_X1 FILLER_81_782 ();
 FILLCELL_X1 FILLER_81_810 ();
 FILLCELL_X1 FILLER_81_835 ();
 FILLCELL_X1 FILLER_81_850 ();
 FILLCELL_X4 FILLER_81_905 ();
 FILLCELL_X1 FILLER_81_909 ();
 FILLCELL_X16 FILLER_81_913 ();
 FILLCELL_X8 FILLER_81_929 ();
 FILLCELL_X1 FILLER_81_937 ();
 FILLCELL_X1 FILLER_81_955 ();
 FILLCELL_X2 FILLER_81_1010 ();
 FILLCELL_X1 FILLER_81_1029 ();
 FILLCELL_X2 FILLER_81_1039 ();
 FILLCELL_X1 FILLER_82_23 ();
 FILLCELL_X4 FILLER_82_56 ();
 FILLCELL_X2 FILLER_82_60 ();
 FILLCELL_X1 FILLER_82_62 ();
 FILLCELL_X2 FILLER_82_70 ();
 FILLCELL_X4 FILLER_82_90 ();
 FILLCELL_X2 FILLER_82_94 ();
 FILLCELL_X1 FILLER_82_100 ();
 FILLCELL_X4 FILLER_82_125 ();
 FILLCELL_X1 FILLER_82_129 ();
 FILLCELL_X8 FILLER_82_146 ();
 FILLCELL_X1 FILLER_82_154 ();
 FILLCELL_X2 FILLER_82_173 ();
 FILLCELL_X2 FILLER_82_216 ();
 FILLCELL_X2 FILLER_82_228 ();
 FILLCELL_X4 FILLER_82_232 ();
 FILLCELL_X4 FILLER_82_276 ();
 FILLCELL_X8 FILLER_82_340 ();
 FILLCELL_X2 FILLER_82_348 ();
 FILLCELL_X16 FILLER_82_370 ();
 FILLCELL_X4 FILLER_82_386 ();
 FILLCELL_X2 FILLER_82_390 ();
 FILLCELL_X1 FILLER_82_479 ();
 FILLCELL_X1 FILLER_82_514 ();
 FILLCELL_X1 FILLER_82_570 ();
 FILLCELL_X2 FILLER_82_595 ();
 FILLCELL_X1 FILLER_82_597 ();
 FILLCELL_X1 FILLER_82_627 ();
 FILLCELL_X1 FILLER_82_639 ();
 FILLCELL_X8 FILLER_82_642 ();
 FILLCELL_X1 FILLER_82_650 ();
 FILLCELL_X4 FILLER_82_659 ();
 FILLCELL_X2 FILLER_82_663 ();
 FILLCELL_X16 FILLER_82_685 ();
 FILLCELL_X2 FILLER_82_701 ();
 FILLCELL_X1 FILLER_82_703 ();
 FILLCELL_X1 FILLER_82_799 ();
 FILLCELL_X1 FILLER_82_840 ();
 FILLCELL_X4 FILLER_82_859 ();
 FILLCELL_X1 FILLER_82_863 ();
 FILLCELL_X4 FILLER_82_878 ();
 FILLCELL_X1 FILLER_82_955 ();
 FILLCELL_X2 FILLER_82_1054 ();
 FILLCELL_X2 FILLER_82_1146 ();
 FILLCELL_X2 FILLER_83_34 ();
 FILLCELL_X4 FILLER_83_51 ();
 FILLCELL_X1 FILLER_83_55 ();
 FILLCELL_X4 FILLER_83_108 ();
 FILLCELL_X2 FILLER_83_112 ();
 FILLCELL_X4 FILLER_83_134 ();
 FILLCELL_X4 FILLER_83_154 ();
 FILLCELL_X1 FILLER_83_158 ();
 FILLCELL_X1 FILLER_83_163 ();
 FILLCELL_X2 FILLER_83_176 ();
 FILLCELL_X2 FILLER_83_180 ();
 FILLCELL_X1 FILLER_83_182 ();
 FILLCELL_X4 FILLER_83_185 ();
 FILLCELL_X2 FILLER_83_189 ();
 FILLCELL_X1 FILLER_83_193 ();
 FILLCELL_X4 FILLER_83_219 ();
 FILLCELL_X2 FILLER_83_223 ();
 FILLCELL_X1 FILLER_83_225 ();
 FILLCELL_X8 FILLER_83_255 ();
 FILLCELL_X2 FILLER_83_263 ();
 FILLCELL_X1 FILLER_83_265 ();
 FILLCELL_X1 FILLER_83_324 ();
 FILLCELL_X8 FILLER_83_371 ();
 FILLCELL_X2 FILLER_83_379 ();
 FILLCELL_X1 FILLER_83_381 ();
 FILLCELL_X1 FILLER_83_521 ();
 FILLCELL_X1 FILLER_83_529 ();
 FILLCELL_X1 FILLER_83_536 ();
 FILLCELL_X1 FILLER_83_554 ();
 FILLCELL_X1 FILLER_83_557 ();
 FILLCELL_X1 FILLER_83_562 ();
 FILLCELL_X1 FILLER_83_565 ();
 FILLCELL_X1 FILLER_83_568 ();
 FILLCELL_X1 FILLER_83_579 ();
 FILLCELL_X2 FILLER_83_618 ();
 FILLCELL_X8 FILLER_83_640 ();
 FILLCELL_X2 FILLER_83_648 ();
 FILLCELL_X2 FILLER_83_670 ();
 FILLCELL_X2 FILLER_83_685 ();
 FILLCELL_X8 FILLER_83_707 ();
 FILLCELL_X1 FILLER_83_715 ();
 FILLCELL_X1 FILLER_83_753 ();
 FILLCELL_X1 FILLER_83_842 ();
 FILLCELL_X1 FILLER_83_853 ();
 FILLCELL_X1 FILLER_83_858 ();
 FILLCELL_X2 FILLER_83_861 ();
 FILLCELL_X16 FILLER_83_875 ();
 FILLCELL_X4 FILLER_83_906 ();
 FILLCELL_X2 FILLER_83_910 ();
 FILLCELL_X2 FILLER_83_936 ();
 FILLCELL_X1 FILLER_83_978 ();
 FILLCELL_X1 FILLER_83_1043 ();
 FILLCELL_X2 FILLER_83_1055 ();
 FILLCELL_X1 FILLER_83_1070 ();
 FILLCELL_X2 FILLER_83_1124 ();
 FILLCELL_X4 FILLER_84_4 ();
 FILLCELL_X8 FILLER_84_73 ();
 FILLCELL_X4 FILLER_84_85 ();
 FILLCELL_X2 FILLER_84_89 ();
 FILLCELL_X4 FILLER_84_93 ();
 FILLCELL_X2 FILLER_84_99 ();
 FILLCELL_X1 FILLER_84_101 ();
 FILLCELL_X2 FILLER_84_110 ();
 FILLCELL_X1 FILLER_84_112 ();
 FILLCELL_X4 FILLER_84_117 ();
 FILLCELL_X1 FILLER_84_121 ();
 FILLCELL_X1 FILLER_84_140 ();
 FILLCELL_X8 FILLER_84_254 ();
 FILLCELL_X1 FILLER_84_262 ();
 FILLCELL_X4 FILLER_84_305 ();
 FILLCELL_X1 FILLER_84_309 ();
 FILLCELL_X2 FILLER_84_330 ();
 FILLCELL_X8 FILLER_84_336 ();
 FILLCELL_X1 FILLER_84_344 ();
 FILLCELL_X16 FILLER_84_367 ();
 FILLCELL_X4 FILLER_84_383 ();
 FILLCELL_X1 FILLER_84_429 ();
 FILLCELL_X1 FILLER_84_501 ();
 FILLCELL_X1 FILLER_84_539 ();
 FILLCELL_X2 FILLER_84_547 ();
 FILLCELL_X1 FILLER_84_605 ();
 FILLCELL_X1 FILLER_84_609 ();
 FILLCELL_X8 FILLER_84_636 ();
 FILLCELL_X4 FILLER_84_664 ();
 FILLCELL_X1 FILLER_84_668 ();
 FILLCELL_X1 FILLER_84_679 ();
 FILLCELL_X2 FILLER_84_715 ();
 FILLCELL_X1 FILLER_84_717 ();
 FILLCELL_X1 FILLER_84_772 ();
 FILLCELL_X2 FILLER_84_821 ();
 FILLCELL_X1 FILLER_84_823 ();
 FILLCELL_X2 FILLER_84_863 ();
 FILLCELL_X8 FILLER_84_885 ();
 FILLCELL_X2 FILLER_84_893 ();
 FILLCELL_X1 FILLER_84_895 ();
 FILLCELL_X2 FILLER_84_999 ();
 FILLCELL_X1 FILLER_84_1001 ();
 FILLCELL_X1 FILLER_84_1016 ();
 FILLCELL_X1 FILLER_84_1024 ();
 FILLCELL_X1 FILLER_84_1032 ();
 FILLCELL_X1 FILLER_84_1055 ();
 FILLCELL_X8 FILLER_84_1106 ();
 FILLCELL_X4 FILLER_84_1114 ();
 FILLCELL_X1 FILLER_84_1118 ();
 FILLCELL_X1 FILLER_85_30 ();
 FILLCELL_X1 FILLER_85_40 ();
 FILLCELL_X2 FILLER_85_45 ();
 FILLCELL_X4 FILLER_85_65 ();
 FILLCELL_X2 FILLER_85_69 ();
 FILLCELL_X4 FILLER_85_73 ();
 FILLCELL_X2 FILLER_85_85 ();
 FILLCELL_X1 FILLER_85_87 ();
 FILLCELL_X4 FILLER_85_122 ();
 FILLCELL_X2 FILLER_85_126 ();
 FILLCELL_X1 FILLER_85_128 ();
 FILLCELL_X1 FILLER_85_133 ();
 FILLCELL_X8 FILLER_85_140 ();
 FILLCELL_X1 FILLER_85_152 ();
 FILLCELL_X1 FILLER_85_160 ();
 FILLCELL_X4 FILLER_85_167 ();
 FILLCELL_X1 FILLER_85_171 ();
 FILLCELL_X4 FILLER_85_190 ();
 FILLCELL_X1 FILLER_85_194 ();
 FILLCELL_X1 FILLER_85_199 ();
 FILLCELL_X2 FILLER_85_202 ();
 FILLCELL_X4 FILLER_85_224 ();
 FILLCELL_X4 FILLER_85_255 ();
 FILLCELL_X2 FILLER_85_259 ();
 FILLCELL_X1 FILLER_85_261 ();
 FILLCELL_X1 FILLER_85_298 ();
 FILLCELL_X2 FILLER_85_311 ();
 FILLCELL_X1 FILLER_85_319 ();
 FILLCELL_X2 FILLER_85_324 ();
 FILLCELL_X1 FILLER_85_326 ();
 FILLCELL_X2 FILLER_85_331 ();
 FILLCELL_X1 FILLER_85_333 ();
 FILLCELL_X4 FILLER_85_356 ();
 FILLCELL_X4 FILLER_85_374 ();
 FILLCELL_X2 FILLER_85_378 ();
 FILLCELL_X1 FILLER_85_511 ();
 FILLCELL_X1 FILLER_85_517 ();
 FILLCELL_X4 FILLER_85_526 ();
 FILLCELL_X2 FILLER_85_530 ();
 FILLCELL_X1 FILLER_85_532 ();
 FILLCELL_X1 FILLER_85_542 ();
 FILLCELL_X1 FILLER_85_547 ();
 FILLCELL_X1 FILLER_85_552 ();
 FILLCELL_X2 FILLER_85_565 ();
 FILLCELL_X1 FILLER_85_574 ();
 FILLCELL_X4 FILLER_85_581 ();
 FILLCELL_X2 FILLER_85_585 ();
 FILLCELL_X2 FILLER_85_616 ();
 FILLCELL_X1 FILLER_85_618 ();
 FILLCELL_X2 FILLER_85_631 ();
 FILLCELL_X1 FILLER_85_633 ();
 FILLCELL_X4 FILLER_85_642 ();
 FILLCELL_X2 FILLER_85_646 ();
 FILLCELL_X1 FILLER_85_648 ();
 FILLCELL_X2 FILLER_85_669 ();
 FILLCELL_X2 FILLER_85_700 ();
 FILLCELL_X1 FILLER_85_702 ();
 FILLCELL_X2 FILLER_85_779 ();
 FILLCELL_X2 FILLER_85_805 ();
 FILLCELL_X4 FILLER_85_827 ();
 FILLCELL_X1 FILLER_85_831 ();
 FILLCELL_X1 FILLER_85_836 ();
 FILLCELL_X4 FILLER_85_839 ();
 FILLCELL_X2 FILLER_85_851 ();
 FILLCELL_X1 FILLER_85_853 ();
 FILLCELL_X2 FILLER_85_872 ();
 FILLCELL_X1 FILLER_85_874 ();
 FILLCELL_X2 FILLER_85_897 ();
 FILLCELL_X1 FILLER_85_921 ();
 FILLCELL_X4 FILLER_85_1085 ();
 FILLCELL_X1 FILLER_85_1089 ();
 FILLCELL_X1 FILLER_85_1141 ();
 FILLCELL_X2 FILLER_85_1145 ();
 FILLCELL_X1 FILLER_85_1147 ();
 FILLCELL_X2 FILLER_86_10 ();
 FILLCELL_X1 FILLER_86_12 ();
 FILLCELL_X1 FILLER_86_50 ();
 FILLCELL_X2 FILLER_86_55 ();
 FILLCELL_X1 FILLER_86_93 ();
 FILLCELL_X4 FILLER_86_97 ();
 FILLCELL_X2 FILLER_86_101 ();
 FILLCELL_X1 FILLER_86_106 ();
 FILLCELL_X2 FILLER_86_110 ();
 FILLCELL_X1 FILLER_86_128 ();
 FILLCELL_X4 FILLER_86_153 ();
 FILLCELL_X2 FILLER_86_157 ();
 FILLCELL_X1 FILLER_86_175 ();
 FILLCELL_X1 FILLER_86_194 ();
 FILLCELL_X1 FILLER_86_254 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X2 FILLER_86_289 ();
 FILLCELL_X1 FILLER_86_319 ();
 FILLCELL_X1 FILLER_86_340 ();
 FILLCELL_X1 FILLER_86_365 ();
 FILLCELL_X2 FILLER_86_371 ();
 FILLCELL_X1 FILLER_86_384 ();
 FILLCELL_X1 FILLER_86_405 ();
 FILLCELL_X1 FILLER_86_423 ();
 FILLCELL_X1 FILLER_86_441 ();
 FILLCELL_X2 FILLER_86_503 ();
 FILLCELL_X2 FILLER_86_569 ();
 FILLCELL_X2 FILLER_86_594 ();
 FILLCELL_X4 FILLER_86_620 ();
 FILLCELL_X1 FILLER_86_632 ();
 FILLCELL_X1 FILLER_86_640 ();
 FILLCELL_X2 FILLER_86_644 ();
 FILLCELL_X1 FILLER_86_676 ();
 FILLCELL_X1 FILLER_86_687 ();
 FILLCELL_X2 FILLER_86_762 ();
 FILLCELL_X1 FILLER_86_771 ();
 FILLCELL_X2 FILLER_86_796 ();
 FILLCELL_X1 FILLER_86_798 ();
 FILLCELL_X4 FILLER_86_828 ();
 FILLCELL_X1 FILLER_86_832 ();
 FILLCELL_X1 FILLER_86_839 ();
 FILLCELL_X4 FILLER_86_858 ();
 FILLCELL_X2 FILLER_86_862 ();
 FILLCELL_X1 FILLER_86_868 ();
 FILLCELL_X8 FILLER_86_889 ();
 FILLCELL_X1 FILLER_86_897 ();
 FILLCELL_X2 FILLER_86_939 ();
 FILLCELL_X1 FILLER_86_956 ();
 FILLCELL_X1 FILLER_86_1057 ();
 FILLCELL_X1 FILLER_86_1065 ();
 FILLCELL_X1 FILLER_86_1083 ();
 FILLCELL_X1 FILLER_86_1110 ();
 FILLCELL_X1 FILLER_87_15 ();
 FILLCELL_X1 FILLER_87_35 ();
 FILLCELL_X1 FILLER_87_38 ();
 FILLCELL_X2 FILLER_87_41 ();
 FILLCELL_X1 FILLER_87_59 ();
 FILLCELL_X4 FILLER_87_111 ();
 FILLCELL_X1 FILLER_87_115 ();
 FILLCELL_X2 FILLER_87_118 ();
 FILLCELL_X4 FILLER_87_124 ();
 FILLCELL_X1 FILLER_87_128 ();
 FILLCELL_X4 FILLER_87_137 ();
 FILLCELL_X2 FILLER_87_141 ();
 FILLCELL_X4 FILLER_87_157 ();
 FILLCELL_X1 FILLER_87_163 ();
 FILLCELL_X1 FILLER_87_168 ();
 FILLCELL_X1 FILLER_87_173 ();
 FILLCELL_X2 FILLER_87_206 ();
 FILLCELL_X1 FILLER_87_208 ();
 FILLCELL_X4 FILLER_87_285 ();
 FILLCELL_X4 FILLER_87_298 ();
 FILLCELL_X2 FILLER_87_302 ();
 FILLCELL_X2 FILLER_87_310 ();
 FILLCELL_X1 FILLER_87_340 ();
 FILLCELL_X1 FILLER_87_363 ();
 FILLCELL_X1 FILLER_87_368 ();
 FILLCELL_X1 FILLER_87_393 ();
 FILLCELL_X1 FILLER_87_414 ();
 FILLCELL_X1 FILLER_87_432 ();
 FILLCELL_X1 FILLER_87_474 ();
 FILLCELL_X1 FILLER_87_491 ();
 FILLCELL_X2 FILLER_87_512 ();
 FILLCELL_X1 FILLER_87_549 ();
 FILLCELL_X1 FILLER_87_554 ();
 FILLCELL_X4 FILLER_87_561 ();
 FILLCELL_X2 FILLER_87_565 ();
 FILLCELL_X1 FILLER_87_578 ();
 FILLCELL_X2 FILLER_87_583 ();
 FILLCELL_X1 FILLER_87_585 ();
 FILLCELL_X1 FILLER_87_603 ();
 FILLCELL_X2 FILLER_87_634 ();
 FILLCELL_X2 FILLER_87_648 ();
 FILLCELL_X4 FILLER_87_670 ();
 FILLCELL_X2 FILLER_87_674 ();
 FILLCELL_X2 FILLER_87_682 ();
 FILLCELL_X1 FILLER_87_687 ();
 FILLCELL_X1 FILLER_87_715 ();
 FILLCELL_X1 FILLER_87_749 ();
 FILLCELL_X1 FILLER_87_820 ();
 FILLCELL_X2 FILLER_87_845 ();
 FILLCELL_X2 FILLER_87_863 ();
 FILLCELL_X1 FILLER_87_867 ();
 FILLCELL_X4 FILLER_87_880 ();
 FILLCELL_X8 FILLER_87_909 ();
 FILLCELL_X1 FILLER_87_917 ();
 FILLCELL_X2 FILLER_87_920 ();
 FILLCELL_X1 FILLER_87_947 ();
 FILLCELL_X1 FILLER_87_952 ();
 FILLCELL_X2 FILLER_87_1033 ();
 FILLCELL_X1 FILLER_87_1121 ();
 FILLCELL_X4 FILLER_88_27 ();
 FILLCELL_X2 FILLER_88_31 ();
 FILLCELL_X1 FILLER_88_33 ();
 FILLCELL_X4 FILLER_88_37 ();
 FILLCELL_X2 FILLER_88_41 ();
 FILLCELL_X2 FILLER_88_45 ();
 FILLCELL_X2 FILLER_88_60 ();
 FILLCELL_X1 FILLER_88_62 ();
 FILLCELL_X2 FILLER_88_65 ();
 FILLCELL_X2 FILLER_88_87 ();
 FILLCELL_X4 FILLER_88_93 ();
 FILLCELL_X2 FILLER_88_97 ();
 FILLCELL_X1 FILLER_88_99 ();
 FILLCELL_X1 FILLER_88_102 ();
 FILLCELL_X1 FILLER_88_139 ();
 FILLCELL_X1 FILLER_88_144 ();
 FILLCELL_X1 FILLER_88_177 ();
 FILLCELL_X2 FILLER_88_188 ();
 FILLCELL_X4 FILLER_88_244 ();
 FILLCELL_X2 FILLER_88_268 ();
 FILLCELL_X1 FILLER_88_270 ();
 FILLCELL_X4 FILLER_88_291 ();
 FILLCELL_X1 FILLER_88_295 ();
 FILLCELL_X1 FILLER_88_322 ();
 FILLCELL_X1 FILLER_88_341 ();
 FILLCELL_X2 FILLER_88_347 ();
 FILLCELL_X1 FILLER_88_349 ();
 FILLCELL_X1 FILLER_88_370 ();
 FILLCELL_X1 FILLER_88_389 ();
 FILLCELL_X1 FILLER_88_401 ();
 FILLCELL_X1 FILLER_88_408 ();
 FILLCELL_X2 FILLER_88_429 ();
 FILLCELL_X1 FILLER_88_431 ();
 FILLCELL_X1 FILLER_88_478 ();
 FILLCELL_X2 FILLER_88_490 ();
 FILLCELL_X2 FILLER_88_514 ();
 FILLCELL_X2 FILLER_88_520 ();
 FILLCELL_X1 FILLER_88_522 ();
 FILLCELL_X1 FILLER_88_545 ();
 FILLCELL_X1 FILLER_88_552 ();
 FILLCELL_X1 FILLER_88_589 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X1 FILLER_88_632 ();
 FILLCELL_X8 FILLER_88_644 ();
 FILLCELL_X1 FILLER_88_672 ();
 FILLCELL_X1 FILLER_88_683 ();
 FILLCELL_X4 FILLER_88_760 ();
 FILLCELL_X1 FILLER_88_778 ();
 FILLCELL_X2 FILLER_88_789 ();
 FILLCELL_X1 FILLER_88_791 ();
 FILLCELL_X4 FILLER_88_826 ();
 FILLCELL_X1 FILLER_88_882 ();
 FILLCELL_X4 FILLER_88_889 ();
 FILLCELL_X2 FILLER_88_893 ();
 FILLCELL_X4 FILLER_88_915 ();
 FILLCELL_X8 FILLER_88_939 ();
 FILLCELL_X1 FILLER_88_1011 ();
 FILLCELL_X1 FILLER_88_1063 ();
 FILLCELL_X4 FILLER_89_42 ();
 FILLCELL_X4 FILLER_89_116 ();
 FILLCELL_X1 FILLER_89_124 ();
 FILLCELL_X1 FILLER_89_145 ();
 FILLCELL_X2 FILLER_89_174 ();
 FILLCELL_X1 FILLER_89_176 ();
 FILLCELL_X32 FILLER_89_200 ();
 FILLCELL_X2 FILLER_89_236 ();
 FILLCELL_X1 FILLER_89_258 ();
 FILLCELL_X2 FILLER_89_300 ();
 FILLCELL_X1 FILLER_89_302 ();
 FILLCELL_X1 FILLER_89_329 ();
 FILLCELL_X1 FILLER_89_354 ();
 FILLCELL_X2 FILLER_89_393 ();
 FILLCELL_X4 FILLER_89_415 ();
 FILLCELL_X1 FILLER_89_419 ();
 FILLCELL_X1 FILLER_89_474 ();
 FILLCELL_X1 FILLER_89_536 ();
 FILLCELL_X1 FILLER_89_584 ();
 FILLCELL_X1 FILLER_89_604 ();
 FILLCELL_X4 FILLER_89_630 ();
 FILLCELL_X2 FILLER_89_634 ();
 FILLCELL_X1 FILLER_89_636 ();
 FILLCELL_X1 FILLER_89_694 ();
 FILLCELL_X1 FILLER_89_752 ();
 FILLCELL_X1 FILLER_89_767 ();
 FILLCELL_X1 FILLER_89_779 ();
 FILLCELL_X2 FILLER_89_784 ();
 FILLCELL_X2 FILLER_89_806 ();
 FILLCELL_X2 FILLER_89_848 ();
 FILLCELL_X1 FILLER_89_855 ();
 FILLCELL_X2 FILLER_89_872 ();
 FILLCELL_X1 FILLER_89_874 ();
 FILLCELL_X2 FILLER_89_881 ();
 FILLCELL_X2 FILLER_89_903 ();
 FILLCELL_X1 FILLER_89_905 ();
 FILLCELL_X2 FILLER_89_926 ();
 FILLCELL_X1 FILLER_89_928 ();
 FILLCELL_X2 FILLER_89_933 ();
 FILLCELL_X2 FILLER_89_949 ();
 FILLCELL_X2 FILLER_89_956 ();
 FILLCELL_X1 FILLER_89_967 ();
 FILLCELL_X1 FILLER_89_989 ();
 FILLCELL_X1 FILLER_89_994 ();
 FILLCELL_X1 FILLER_89_1077 ();
 FILLCELL_X1 FILLER_89_1132 ();
 FILLCELL_X8 FILLER_89_1140 ();
 FILLCELL_X1 FILLER_90_23 ();
 FILLCELL_X2 FILLER_90_28 ();
 FILLCELL_X4 FILLER_90_56 ();
 FILLCELL_X2 FILLER_90_60 ();
 FILLCELL_X1 FILLER_90_65 ();
 FILLCELL_X2 FILLER_90_93 ();
 FILLCELL_X4 FILLER_90_97 ();
 FILLCELL_X2 FILLER_90_101 ();
 FILLCELL_X8 FILLER_90_105 ();
 FILLCELL_X2 FILLER_90_113 ();
 FILLCELL_X1 FILLER_90_115 ();
 FILLCELL_X1 FILLER_90_165 ();
 FILLCELL_X1 FILLER_90_170 ();
 FILLCELL_X1 FILLER_90_183 ();
 FILLCELL_X2 FILLER_90_187 ();
 FILLCELL_X1 FILLER_90_189 ();
 FILLCELL_X4 FILLER_90_198 ();
 FILLCELL_X2 FILLER_90_204 ();
 FILLCELL_X4 FILLER_90_208 ();
 FILLCELL_X1 FILLER_90_212 ();
 FILLCELL_X2 FILLER_90_283 ();
 FILLCELL_X4 FILLER_90_287 ();
 FILLCELL_X2 FILLER_90_291 ();
 FILLCELL_X1 FILLER_90_300 ();
 FILLCELL_X1 FILLER_90_308 ();
 FILLCELL_X1 FILLER_90_313 ();
 FILLCELL_X1 FILLER_90_321 ();
 FILLCELL_X1 FILLER_90_349 ();
 FILLCELL_X2 FILLER_90_353 ();
 FILLCELL_X2 FILLER_90_411 ();
 FILLCELL_X32 FILLER_90_421 ();
 FILLCELL_X4 FILLER_90_453 ();
 FILLCELL_X4 FILLER_90_499 ();
 FILLCELL_X2 FILLER_90_503 ();
 FILLCELL_X1 FILLER_90_513 ();
 FILLCELL_X1 FILLER_90_558 ();
 FILLCELL_X1 FILLER_90_566 ();
 FILLCELL_X1 FILLER_90_576 ();
 FILLCELL_X1 FILLER_90_587 ();
 FILLCELL_X1 FILLER_90_608 ();
 FILLCELL_X2 FILLER_90_676 ();
 FILLCELL_X2 FILLER_90_686 ();
 FILLCELL_X1 FILLER_90_688 ();
 FILLCELL_X2 FILLER_90_734 ();
 FILLCELL_X1 FILLER_90_817 ();
 FILLCELL_X8 FILLER_90_864 ();
 FILLCELL_X4 FILLER_90_872 ();
 FILLCELL_X2 FILLER_90_876 ();
 FILLCELL_X1 FILLER_90_940 ();
 FILLCELL_X2 FILLER_90_1001 ();
 FILLCELL_X1 FILLER_90_1043 ();
 FILLCELL_X2 FILLER_90_1065 ();
 FILLCELL_X1 FILLER_90_1103 ();
 FILLCELL_X2 FILLER_90_1138 ();
 FILLCELL_X4 FILLER_90_1144 ();
 FILLCELL_X1 FILLER_91_22 ();
 FILLCELL_X1 FILLER_91_41 ();
 FILLCELL_X8 FILLER_91_88 ();
 FILLCELL_X2 FILLER_91_96 ();
 FILLCELL_X2 FILLER_91_118 ();
 FILLCELL_X1 FILLER_91_120 ();
 FILLCELL_X2 FILLER_91_135 ();
 FILLCELL_X1 FILLER_91_171 ();
 FILLCELL_X4 FILLER_91_181 ();
 FILLCELL_X2 FILLER_91_185 ();
 FILLCELL_X2 FILLER_91_247 ();
 FILLCELL_X1 FILLER_91_262 ();
 FILLCELL_X2 FILLER_91_273 ();
 FILLCELL_X4 FILLER_91_281 ();
 FILLCELL_X1 FILLER_91_285 ();
 FILLCELL_X2 FILLER_91_368 ();
 FILLCELL_X1 FILLER_91_374 ();
 FILLCELL_X1 FILLER_91_383 ();
 FILLCELL_X2 FILLER_91_388 ();
 FILLCELL_X1 FILLER_91_390 ();
 FILLCELL_X4 FILLER_91_462 ();
 FILLCELL_X2 FILLER_91_470 ();
 FILLCELL_X1 FILLER_91_498 ();
 FILLCELL_X1 FILLER_91_534 ();
 FILLCELL_X4 FILLER_91_588 ();
 FILLCELL_X4 FILLER_91_634 ();
 FILLCELL_X2 FILLER_91_638 ();
 FILLCELL_X1 FILLER_91_670 ();
 FILLCELL_X1 FILLER_91_673 ();
 FILLCELL_X1 FILLER_91_684 ();
 FILLCELL_X1 FILLER_91_798 ();
 FILLCELL_X1 FILLER_91_803 ();
 FILLCELL_X1 FILLER_91_806 ();
 FILLCELL_X1 FILLER_91_809 ();
 FILLCELL_X1 FILLER_91_816 ();
 FILLCELL_X1 FILLER_91_826 ();
 FILLCELL_X8 FILLER_91_851 ();
 FILLCELL_X2 FILLER_91_859 ();
 FILLCELL_X16 FILLER_91_864 ();
 FILLCELL_X8 FILLER_91_880 ();
 FILLCELL_X2 FILLER_91_888 ();
 FILLCELL_X16 FILLER_91_910 ();
 FILLCELL_X4 FILLER_91_926 ();
 FILLCELL_X2 FILLER_91_930 ();
 FILLCELL_X1 FILLER_91_951 ();
 FILLCELL_X1 FILLER_91_959 ();
 FILLCELL_X1 FILLER_91_967 ();
 FILLCELL_X1 FILLER_91_980 ();
 FILLCELL_X1 FILLER_91_1007 ();
 FILLCELL_X1 FILLER_91_1015 ();
 FILLCELL_X1 FILLER_91_1023 ();
 FILLCELL_X2 FILLER_91_1061 ();
 FILLCELL_X2 FILLER_91_1105 ();
 FILLCELL_X2 FILLER_91_1116 ();
 FILLCELL_X1 FILLER_91_1118 ();
 FILLCELL_X1 FILLER_91_1124 ();
 FILLCELL_X4 FILLER_91_1144 ();
 FILLCELL_X2 FILLER_92_1 ();
 FILLCELL_X1 FILLER_92_3 ();
 FILLCELL_X1 FILLER_92_6 ();
 FILLCELL_X2 FILLER_92_23 ();
 FILLCELL_X1 FILLER_92_25 ();
 FILLCELL_X2 FILLER_92_28 ();
 FILLCELL_X4 FILLER_92_54 ();
 FILLCELL_X2 FILLER_92_58 ();
 FILLCELL_X4 FILLER_92_62 ();
 FILLCELL_X2 FILLER_92_66 ();
 FILLCELL_X1 FILLER_92_68 ();
 FILLCELL_X2 FILLER_92_133 ();
 FILLCELL_X1 FILLER_92_135 ();
 FILLCELL_X4 FILLER_92_185 ();
 FILLCELL_X2 FILLER_92_193 ();
 FILLCELL_X4 FILLER_92_215 ();
 FILLCELL_X1 FILLER_92_229 ();
 FILLCELL_X1 FILLER_92_237 ();
 FILLCELL_X2 FILLER_92_260 ();
 FILLCELL_X2 FILLER_92_389 ();
 FILLCELL_X2 FILLER_92_402 ();
 FILLCELL_X1 FILLER_92_417 ();
 FILLCELL_X1 FILLER_92_453 ();
 FILLCELL_X1 FILLER_92_461 ();
 FILLCELL_X2 FILLER_92_466 ();
 FILLCELL_X1 FILLER_92_475 ();
 FILLCELL_X4 FILLER_92_483 ();
 FILLCELL_X2 FILLER_92_619 ();
 FILLCELL_X1 FILLER_92_642 ();
 FILLCELL_X1 FILLER_92_652 ();
 FILLCELL_X2 FILLER_92_658 ();
 FILLCELL_X2 FILLER_92_665 ();
 FILLCELL_X1 FILLER_92_667 ();
 FILLCELL_X2 FILLER_92_671 ();
 FILLCELL_X1 FILLER_92_681 ();
 FILLCELL_X2 FILLER_92_701 ();
 FILLCELL_X1 FILLER_92_703 ();
 FILLCELL_X4 FILLER_92_773 ();
 FILLCELL_X8 FILLER_92_875 ();
 FILLCELL_X4 FILLER_92_908 ();
 FILLCELL_X2 FILLER_92_912 ();
 FILLCELL_X1 FILLER_92_914 ();
 FILLCELL_X1 FILLER_92_955 ();
 FILLCELL_X1 FILLER_92_979 ();
 FILLCELL_X2 FILLER_92_991 ();
 FILLCELL_X1 FILLER_92_1030 ();
 FILLCELL_X1 FILLER_92_1040 ();
 FILLCELL_X2 FILLER_92_1084 ();
 FILLCELL_X1 FILLER_92_1086 ();
 FILLCELL_X1 FILLER_92_1090 ();
 FILLCELL_X4 FILLER_92_1131 ();
 FILLCELL_X8 FILLER_92_1139 ();
 FILLCELL_X1 FILLER_92_1147 ();
 FILLCELL_X1 FILLER_93_1 ();
 FILLCELL_X2 FILLER_93_5 ();
 FILLCELL_X2 FILLER_93_11 ();
 FILLCELL_X16 FILLER_93_77 ();
 FILLCELL_X8 FILLER_93_93 ();
 FILLCELL_X4 FILLER_93_101 ();
 FILLCELL_X2 FILLER_93_105 ();
 FILLCELL_X32 FILLER_93_110 ();
 FILLCELL_X8 FILLER_93_142 ();
 FILLCELL_X4 FILLER_93_150 ();
 FILLCELL_X2 FILLER_93_154 ();
 FILLCELL_X1 FILLER_93_163 ();
 FILLCELL_X1 FILLER_93_176 ();
 FILLCELL_X1 FILLER_93_179 ();
 FILLCELL_X1 FILLER_93_200 ();
 FILLCELL_X1 FILLER_93_221 ();
 FILLCELL_X2 FILLER_93_282 ();
 FILLCELL_X4 FILLER_93_372 ();
 FILLCELL_X1 FILLER_93_392 ();
 FILLCELL_X1 FILLER_93_399 ();
 FILLCELL_X2 FILLER_93_403 ();
 FILLCELL_X1 FILLER_93_405 ();
 FILLCELL_X16 FILLER_93_425 ();
 FILLCELL_X8 FILLER_93_441 ();
 FILLCELL_X2 FILLER_93_449 ();
 FILLCELL_X1 FILLER_93_455 ();
 FILLCELL_X1 FILLER_93_463 ();
 FILLCELL_X1 FILLER_93_471 ();
 FILLCELL_X2 FILLER_93_479 ();
 FILLCELL_X1 FILLER_93_481 ();
 FILLCELL_X1 FILLER_93_556 ();
 FILLCELL_X2 FILLER_93_598 ();
 FILLCELL_X2 FILLER_93_695 ();
 FILLCELL_X1 FILLER_93_701 ();
 FILLCELL_X1 FILLER_93_734 ();
 FILLCELL_X2 FILLER_93_783 ();
 FILLCELL_X1 FILLER_93_854 ();
 FILLCELL_X16 FILLER_93_872 ();
 FILLCELL_X4 FILLER_93_888 ();
 FILLCELL_X1 FILLER_93_892 ();
 FILLCELL_X2 FILLER_93_941 ();
 FILLCELL_X4 FILLER_93_949 ();
 FILLCELL_X2 FILLER_93_953 ();
 FILLCELL_X1 FILLER_93_955 ();
 FILLCELL_X4 FILLER_93_958 ();
 FILLCELL_X2 FILLER_93_962 ();
 FILLCELL_X1 FILLER_93_971 ();
 FILLCELL_X1 FILLER_93_975 ();
 FILLCELL_X1 FILLER_93_979 ();
 FILLCELL_X1 FILLER_93_991 ();
 FILLCELL_X2 FILLER_93_996 ();
 FILLCELL_X2 FILLER_93_1032 ();
 FILLCELL_X2 FILLER_93_1036 ();
 FILLCELL_X1 FILLER_93_1038 ();
 FILLCELL_X1 FILLER_93_1095 ();
 FILLCELL_X2 FILLER_93_1100 ();
 FILLCELL_X4 FILLER_93_1127 ();
 FILLCELL_X2 FILLER_93_1131 ();
 FILLCELL_X1 FILLER_93_1133 ();
 FILLCELL_X8 FILLER_93_1137 ();
 FILLCELL_X2 FILLER_93_1145 ();
 FILLCELL_X1 FILLER_93_1147 ();
 FILLCELL_X4 FILLER_94_1 ();
 FILLCELL_X8 FILLER_94_7 ();
 FILLCELL_X4 FILLER_94_34 ();
 FILLCELL_X2 FILLER_94_40 ();
 FILLCELL_X1 FILLER_94_42 ();
 FILLCELL_X2 FILLER_94_47 ();
 FILLCELL_X4 FILLER_94_69 ();
 FILLCELL_X1 FILLER_94_81 ();
 FILLCELL_X1 FILLER_94_86 ();
 FILLCELL_X1 FILLER_94_111 ();
 FILLCELL_X1 FILLER_94_177 ();
 FILLCELL_X2 FILLER_94_185 ();
 FILLCELL_X1 FILLER_94_187 ();
 FILLCELL_X4 FILLER_94_208 ();
 FILLCELL_X1 FILLER_94_212 ();
 FILLCELL_X1 FILLER_94_229 ();
 FILLCELL_X2 FILLER_94_328 ();
 FILLCELL_X2 FILLER_94_391 ();
 FILLCELL_X2 FILLER_94_407 ();
 FILLCELL_X1 FILLER_94_409 ();
 FILLCELL_X4 FILLER_94_426 ();
 FILLCELL_X1 FILLER_94_489 ();
 FILLCELL_X1 FILLER_94_516 ();
 FILLCELL_X1 FILLER_94_568 ();
 FILLCELL_X1 FILLER_94_572 ();
 FILLCELL_X1 FILLER_94_590 ();
 FILLCELL_X4 FILLER_94_617 ();
 FILLCELL_X2 FILLER_94_719 ();
 FILLCELL_X4 FILLER_94_760 ();
 FILLCELL_X2 FILLER_94_805 ();
 FILLCELL_X4 FILLER_94_878 ();
 FILLCELL_X1 FILLER_94_882 ();
 FILLCELL_X4 FILLER_94_950 ();
 FILLCELL_X2 FILLER_94_954 ();
 FILLCELL_X1 FILLER_94_966 ();
 FILLCELL_X2 FILLER_94_971 ();
 FILLCELL_X2 FILLER_94_1029 ();
 FILLCELL_X2 FILLER_94_1045 ();
 FILLCELL_X1 FILLER_94_1067 ();
 FILLCELL_X1 FILLER_94_1109 ();
 FILLCELL_X4 FILLER_94_1124 ();
 FILLCELL_X2 FILLER_94_1128 ();
 FILLCELL_X1 FILLER_94_1130 ();
 FILLCELL_X2 FILLER_94_1137 ();
 FILLCELL_X1 FILLER_94_1139 ();
 FILLCELL_X4 FILLER_94_1143 ();
 FILLCELL_X1 FILLER_94_1147 ();
 FILLCELL_X2 FILLER_95_19 ();
 FILLCELL_X1 FILLER_95_21 ();
 FILLCELL_X1 FILLER_95_38 ();
 FILLCELL_X2 FILLER_95_55 ();
 FILLCELL_X8 FILLER_95_59 ();
 FILLCELL_X2 FILLER_95_69 ();
 FILLCELL_X1 FILLER_95_87 ();
 FILLCELL_X4 FILLER_95_104 ();
 FILLCELL_X2 FILLER_95_130 ();
 FILLCELL_X1 FILLER_95_132 ();
 FILLCELL_X2 FILLER_95_185 ();
 FILLCELL_X2 FILLER_95_191 ();
 FILLCELL_X1 FILLER_95_193 ();
 FILLCELL_X2 FILLER_95_198 ();
 FILLCELL_X1 FILLER_95_200 ();
 FILLCELL_X2 FILLER_95_221 ();
 FILLCELL_X1 FILLER_95_223 ();
 FILLCELL_X1 FILLER_95_229 ();
 FILLCELL_X1 FILLER_95_250 ();
 FILLCELL_X1 FILLER_95_327 ();
 FILLCELL_X1 FILLER_95_368 ();
 FILLCELL_X2 FILLER_95_399 ();
 FILLCELL_X1 FILLER_95_404 ();
 FILLCELL_X8 FILLER_95_412 ();
 FILLCELL_X4 FILLER_95_420 ();
 FILLCELL_X2 FILLER_95_424 ();
 FILLCELL_X1 FILLER_95_459 ();
 FILLCELL_X1 FILLER_95_464 ();
 FILLCELL_X1 FILLER_95_472 ();
 FILLCELL_X1 FILLER_95_507 ();
 FILLCELL_X1 FILLER_95_575 ();
 FILLCELL_X1 FILLER_95_581 ();
 FILLCELL_X1 FILLER_95_602 ();
 FILLCELL_X1 FILLER_95_605 ();
 FILLCELL_X1 FILLER_95_617 ();
 FILLCELL_X1 FILLER_95_631 ();
 FILLCELL_X1 FILLER_95_642 ();
 FILLCELL_X2 FILLER_95_648 ();
 FILLCELL_X1 FILLER_95_672 ();
 FILLCELL_X1 FILLER_95_698 ();
 FILLCELL_X1 FILLER_95_834 ();
 FILLCELL_X2 FILLER_95_877 ();
 FILLCELL_X2 FILLER_95_923 ();
 FILLCELL_X8 FILLER_95_937 ();
 FILLCELL_X1 FILLER_95_945 ();
 FILLCELL_X2 FILLER_95_1034 ();
 FILLCELL_X1 FILLER_95_1036 ();
 FILLCELL_X1 FILLER_95_1054 ();
 FILLCELL_X4 FILLER_95_1058 ();
 FILLCELL_X2 FILLER_95_1062 ();
 FILLCELL_X8 FILLER_95_1095 ();
 FILLCELL_X2 FILLER_95_1103 ();
 FILLCELL_X1 FILLER_95_1105 ();
 FILLCELL_X32 FILLER_95_1109 ();
 FILLCELL_X4 FILLER_95_1141 ();
 FILLCELL_X2 FILLER_95_1145 ();
 FILLCELL_X1 FILLER_95_1147 ();
 FILLCELL_X1 FILLER_96_1 ();
 FILLCELL_X8 FILLER_96_24 ();
 FILLCELL_X8 FILLER_96_34 ();
 FILLCELL_X2 FILLER_96_42 ();
 FILLCELL_X1 FILLER_96_44 ();
 FILLCELL_X2 FILLER_96_49 ();
 FILLCELL_X1 FILLER_96_51 ();
 FILLCELL_X8 FILLER_96_86 ();
 FILLCELL_X16 FILLER_96_116 ();
 FILLCELL_X1 FILLER_96_132 ();
 FILLCELL_X4 FILLER_96_164 ();
 FILLCELL_X2 FILLER_96_171 ();
 FILLCELL_X1 FILLER_96_173 ();
 FILLCELL_X1 FILLER_96_181 ();
 FILLCELL_X8 FILLER_96_192 ();
 FILLCELL_X2 FILLER_96_200 ();
 FILLCELL_X16 FILLER_96_207 ();
 FILLCELL_X1 FILLER_96_223 ();
 FILLCELL_X4 FILLER_96_234 ();
 FILLCELL_X2 FILLER_96_238 ();
 FILLCELL_X1 FILLER_96_260 ();
 FILLCELL_X1 FILLER_96_270 ();
 FILLCELL_X1 FILLER_96_284 ();
 FILLCELL_X2 FILLER_96_299 ();
 FILLCELL_X1 FILLER_96_322 ();
 FILLCELL_X2 FILLER_96_370 ();
 FILLCELL_X1 FILLER_96_390 ();
 FILLCELL_X1 FILLER_96_410 ();
 FILLCELL_X1 FILLER_96_414 ();
 FILLCELL_X1 FILLER_96_427 ();
 FILLCELL_X1 FILLER_96_432 ();
 FILLCELL_X1 FILLER_96_455 ();
 FILLCELL_X1 FILLER_96_463 ();
 FILLCELL_X4 FILLER_96_584 ();
 FILLCELL_X2 FILLER_96_588 ();
 FILLCELL_X1 FILLER_96_590 ();
 FILLCELL_X1 FILLER_96_598 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X1 FILLER_96_702 ();
 FILLCELL_X1 FILLER_96_818 ();
 FILLCELL_X1 FILLER_96_857 ();
 FILLCELL_X1 FILLER_96_883 ();
 FILLCELL_X1 FILLER_96_904 ();
 FILLCELL_X4 FILLER_96_940 ();
 FILLCELL_X1 FILLER_96_946 ();
 FILLCELL_X2 FILLER_96_957 ();
 FILLCELL_X1 FILLER_96_959 ();
 FILLCELL_X2 FILLER_96_964 ();
 FILLCELL_X1 FILLER_96_966 ();
 FILLCELL_X1 FILLER_96_969 ();
 FILLCELL_X2 FILLER_96_978 ();
 FILLCELL_X1 FILLER_96_1066 ();
 FILLCELL_X2 FILLER_96_1071 ();
 FILLCELL_X8 FILLER_96_1086 ();
 FILLCELL_X4 FILLER_96_1094 ();
 FILLCELL_X32 FILLER_96_1104 ();
 FILLCELL_X8 FILLER_96_1136 ();
 FILLCELL_X4 FILLER_96_1144 ();
 FILLCELL_X2 FILLER_97_19 ();
 FILLCELL_X2 FILLER_97_29 ();
 FILLCELL_X1 FILLER_97_31 ();
 FILLCELL_X2 FILLER_97_48 ();
 FILLCELL_X1 FILLER_97_50 ();
 FILLCELL_X4 FILLER_97_63 ();
 FILLCELL_X2 FILLER_97_67 ();
 FILLCELL_X16 FILLER_97_88 ();
 FILLCELL_X2 FILLER_97_106 ();
 FILLCELL_X1 FILLER_97_113 ();
 FILLCELL_X4 FILLER_97_134 ();
 FILLCELL_X2 FILLER_97_138 ();
 FILLCELL_X2 FILLER_97_161 ();
 FILLCELL_X1 FILLER_97_163 ();
 FILLCELL_X1 FILLER_97_194 ();
 FILLCELL_X4 FILLER_97_219 ();
 FILLCELL_X1 FILLER_97_245 ();
 FILLCELL_X2 FILLER_97_276 ();
 FILLCELL_X1 FILLER_97_339 ();
 FILLCELL_X2 FILLER_97_375 ();
 FILLCELL_X1 FILLER_97_396 ();
 FILLCELL_X2 FILLER_97_415 ();
 FILLCELL_X1 FILLER_97_417 ();
 FILLCELL_X1 FILLER_97_434 ();
 FILLCELL_X2 FILLER_97_463 ();
 FILLCELL_X1 FILLER_97_465 ();
 FILLCELL_X1 FILLER_97_570 ();
 FILLCELL_X1 FILLER_97_591 ();
 FILLCELL_X1 FILLER_97_594 ();
 FILLCELL_X1 FILLER_97_609 ();
 FILLCELL_X2 FILLER_97_704 ();
 FILLCELL_X1 FILLER_97_736 ();
 FILLCELL_X2 FILLER_97_812 ();
 FILLCELL_X2 FILLER_97_883 ();
 FILLCELL_X2 FILLER_97_943 ();
 FILLCELL_X1 FILLER_97_995 ();
 FILLCELL_X2 FILLER_97_1074 ();
 FILLCELL_X1 FILLER_97_1076 ();
 FILLCELL_X4 FILLER_97_1084 ();
 FILLCELL_X2 FILLER_97_1088 ();
 FILLCELL_X32 FILLER_97_1114 ();
 FILLCELL_X2 FILLER_97_1146 ();
 FILLCELL_X4 FILLER_98_1 ();
 FILLCELL_X1 FILLER_98_5 ();
 FILLCELL_X4 FILLER_98_41 ();
 FILLCELL_X4 FILLER_98_59 ();
 FILLCELL_X2 FILLER_98_63 ();
 FILLCELL_X1 FILLER_98_81 ();
 FILLCELL_X1 FILLER_98_102 ();
 FILLCELL_X1 FILLER_98_105 ();
 FILLCELL_X4 FILLER_98_126 ();
 FILLCELL_X2 FILLER_98_130 ();
 FILLCELL_X1 FILLER_98_132 ();
 FILLCELL_X2 FILLER_98_143 ();
 FILLCELL_X2 FILLER_98_157 ();
 FILLCELL_X2 FILLER_98_179 ();
 FILLCELL_X1 FILLER_98_195 ();
 FILLCELL_X4 FILLER_98_202 ();
 FILLCELL_X2 FILLER_98_206 ();
 FILLCELL_X8 FILLER_98_228 ();
 FILLCELL_X1 FILLER_98_256 ();
 FILLCELL_X2 FILLER_98_292 ();
 FILLCELL_X1 FILLER_98_336 ();
 FILLCELL_X1 FILLER_98_387 ();
 FILLCELL_X1 FILLER_98_397 ();
 FILLCELL_X2 FILLER_98_401 ();
 FILLCELL_X1 FILLER_98_412 ();
 FILLCELL_X1 FILLER_98_426 ();
 FILLCELL_X1 FILLER_98_430 ();
 FILLCELL_X1 FILLER_98_439 ();
 FILLCELL_X1 FILLER_98_460 ();
 FILLCELL_X2 FILLER_98_528 ();
 FILLCELL_X1 FILLER_98_575 ();
 FILLCELL_X1 FILLER_98_594 ();
 FILLCELL_X1 FILLER_98_632 ();
 FILLCELL_X1 FILLER_98_637 ();
 FILLCELL_X2 FILLER_98_703 ();
 FILLCELL_X1 FILLER_98_846 ();
 FILLCELL_X2 FILLER_98_858 ();
 FILLCELL_X2 FILLER_98_882 ();
 FILLCELL_X1 FILLER_98_903 ();
 FILLCELL_X2 FILLER_98_935 ();
 FILLCELL_X1 FILLER_98_946 ();
 FILLCELL_X1 FILLER_98_953 ();
 FILLCELL_X1 FILLER_98_964 ();
 FILLCELL_X1 FILLER_98_969 ();
 FILLCELL_X1 FILLER_98_974 ();
 FILLCELL_X1 FILLER_98_977 ();
 FILLCELL_X1 FILLER_98_1028 ();
 FILLCELL_X2 FILLER_98_1068 ();
 FILLCELL_X2 FILLER_98_1077 ();
 FILLCELL_X4 FILLER_98_1102 ();
 FILLCELL_X2 FILLER_98_1106 ();
 FILLCELL_X1 FILLER_98_1108 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X4 FILLER_98_1144 ();
 FILLCELL_X1 FILLER_99_1 ();
 FILLCELL_X1 FILLER_99_20 ();
 FILLCELL_X2 FILLER_99_27 ();
 FILLCELL_X1 FILLER_99_29 ();
 FILLCELL_X2 FILLER_99_54 ();
 FILLCELL_X2 FILLER_99_76 ();
 FILLCELL_X1 FILLER_99_78 ();
 FILLCELL_X4 FILLER_99_135 ();
 FILLCELL_X2 FILLER_99_139 ();
 FILLCELL_X2 FILLER_99_149 ();
 FILLCELL_X1 FILLER_99_198 ();
 FILLCELL_X1 FILLER_99_205 ();
 FILLCELL_X4 FILLER_99_212 ();
 FILLCELL_X1 FILLER_99_265 ();
 FILLCELL_X2 FILLER_99_324 ();
 FILLCELL_X1 FILLER_99_379 ();
 FILLCELL_X1 FILLER_99_390 ();
 FILLCELL_X1 FILLER_99_406 ();
 FILLCELL_X1 FILLER_99_424 ();
 FILLCELL_X1 FILLER_99_429 ();
 FILLCELL_X2 FILLER_99_434 ();
 FILLCELL_X4 FILLER_99_458 ();
 FILLCELL_X1 FILLER_99_469 ();
 FILLCELL_X2 FILLER_99_518 ();
 FILLCELL_X2 FILLER_99_566 ();
 FILLCELL_X1 FILLER_99_599 ();
 FILLCELL_X1 FILLER_99_604 ();
 FILLCELL_X4 FILLER_99_627 ();
 FILLCELL_X2 FILLER_99_660 ();
 FILLCELL_X1 FILLER_99_666 ();
 FILLCELL_X2 FILLER_99_671 ();
 FILLCELL_X2 FILLER_99_694 ();
 FILLCELL_X1 FILLER_99_754 ();
 FILLCELL_X1 FILLER_99_868 ();
 FILLCELL_X1 FILLER_99_879 ();
 FILLCELL_X1 FILLER_99_902 ();
 FILLCELL_X2 FILLER_99_920 ();
 FILLCELL_X1 FILLER_99_940 ();
 FILLCELL_X1 FILLER_99_965 ();
 FILLCELL_X1 FILLER_99_1002 ();
 FILLCELL_X1 FILLER_99_1020 ();
 FILLCELL_X2 FILLER_99_1037 ();
 FILLCELL_X1 FILLER_99_1087 ();
 FILLCELL_X1 FILLER_99_1106 ();
 FILLCELL_X32 FILLER_99_1111 ();
 FILLCELL_X4 FILLER_99_1143 ();
 FILLCELL_X1 FILLER_99_1147 ();
 FILLCELL_X4 FILLER_100_1 ();
 FILLCELL_X2 FILLER_100_5 ();
 FILLCELL_X1 FILLER_100_23 ();
 FILLCELL_X1 FILLER_100_44 ();
 FILLCELL_X2 FILLER_100_47 ();
 FILLCELL_X2 FILLER_100_69 ();
 FILLCELL_X1 FILLER_100_105 ();
 FILLCELL_X4 FILLER_100_126 ();
 FILLCELL_X2 FILLER_100_150 ();
 FILLCELL_X1 FILLER_100_152 ();
 FILLCELL_X2 FILLER_100_156 ();
 FILLCELL_X2 FILLER_100_210 ();
 FILLCELL_X4 FILLER_100_226 ();
 FILLCELL_X8 FILLER_100_245 ();
 FILLCELL_X4 FILLER_100_253 ();
 FILLCELL_X1 FILLER_100_257 ();
 FILLCELL_X2 FILLER_100_378 ();
 FILLCELL_X1 FILLER_100_388 ();
 FILLCELL_X1 FILLER_100_409 ();
 FILLCELL_X1 FILLER_100_413 ();
 FILLCELL_X8 FILLER_100_440 ();
 FILLCELL_X2 FILLER_100_448 ();
 FILLCELL_X1 FILLER_100_473 ();
 FILLCELL_X1 FILLER_100_493 ();
 FILLCELL_X1 FILLER_100_576 ();
 FILLCELL_X1 FILLER_100_583 ();
 FILLCELL_X1 FILLER_100_591 ();
 FILLCELL_X2 FILLER_100_598 ();
 FILLCELL_X1 FILLER_100_614 ();
 FILLCELL_X1 FILLER_100_622 ();
 FILLCELL_X1 FILLER_100_630 ();
 FILLCELL_X1 FILLER_100_640 ();
 FILLCELL_X2 FILLER_100_700 ();
 FILLCELL_X2 FILLER_100_768 ();
 FILLCELL_X1 FILLER_100_814 ();
 FILLCELL_X2 FILLER_100_819 ();
 FILLCELL_X1 FILLER_100_821 ();
 FILLCELL_X2 FILLER_100_836 ();
 FILLCELL_X1 FILLER_100_931 ();
 FILLCELL_X1 FILLER_100_993 ();
 FILLCELL_X8 FILLER_100_1028 ();
 FILLCELL_X4 FILLER_100_1036 ();
 FILLCELL_X1 FILLER_100_1040 ();
 FILLCELL_X1 FILLER_100_1061 ();
 FILLCELL_X1 FILLER_100_1086 ();
 FILLCELL_X1 FILLER_100_1094 ();
 FILLCELL_X1 FILLER_100_1098 ();
 FILLCELL_X16 FILLER_100_1122 ();
 FILLCELL_X8 FILLER_100_1138 ();
 FILLCELL_X2 FILLER_100_1146 ();
 FILLCELL_X4 FILLER_101_1 ();
 FILLCELL_X1 FILLER_101_8 ();
 FILLCELL_X2 FILLER_101_19 ();
 FILLCELL_X1 FILLER_101_28 ();
 FILLCELL_X2 FILLER_101_37 ();
 FILLCELL_X1 FILLER_101_39 ();
 FILLCELL_X4 FILLER_101_60 ();
 FILLCELL_X2 FILLER_101_64 ();
 FILLCELL_X1 FILLER_101_66 ();
 FILLCELL_X2 FILLER_101_83 ();
 FILLCELL_X1 FILLER_101_89 ();
 FILLCELL_X4 FILLER_101_108 ();
 FILLCELL_X1 FILLER_101_114 ();
 FILLCELL_X1 FILLER_101_181 ();
 FILLCELL_X1 FILLER_101_188 ();
 FILLCELL_X1 FILLER_101_194 ();
 FILLCELL_X1 FILLER_101_199 ();
 FILLCELL_X4 FILLER_101_208 ();
 FILLCELL_X1 FILLER_101_239 ();
 FILLCELL_X1 FILLER_101_262 ();
 FILLCELL_X1 FILLER_101_357 ();
 FILLCELL_X1 FILLER_101_378 ();
 FILLCELL_X1 FILLER_101_389 ();
 FILLCELL_X1 FILLER_101_394 ();
 FILLCELL_X1 FILLER_101_431 ();
 FILLCELL_X1 FILLER_101_438 ();
 FILLCELL_X1 FILLER_101_449 ();
 FILLCELL_X1 FILLER_101_491 ();
 FILLCELL_X2 FILLER_101_587 ();
 FILLCELL_X1 FILLER_101_589 ();
 FILLCELL_X1 FILLER_101_606 ();
 FILLCELL_X2 FILLER_101_672 ();
 FILLCELL_X1 FILLER_101_678 ();
 FILLCELL_X4 FILLER_101_682 ();
 FILLCELL_X1 FILLER_101_686 ();
 FILLCELL_X1 FILLER_101_711 ();
 FILLCELL_X1 FILLER_101_726 ();
 FILLCELL_X1 FILLER_101_781 ();
 FILLCELL_X1 FILLER_101_802 ();
 FILLCELL_X1 FILLER_101_806 ();
 FILLCELL_X1 FILLER_101_856 ();
 FILLCELL_X1 FILLER_101_894 ();
 FILLCELL_X1 FILLER_101_902 ();
 FILLCELL_X1 FILLER_101_951 ();
 FILLCELL_X2 FILLER_101_954 ();
 FILLCELL_X1 FILLER_101_956 ();
 FILLCELL_X1 FILLER_101_961 ();
 FILLCELL_X1 FILLER_101_1016 ();
 FILLCELL_X1 FILLER_101_1025 ();
 FILLCELL_X2 FILLER_101_1105 ();
 FILLCELL_X2 FILLER_101_1114 ();
 FILLCELL_X16 FILLER_101_1127 ();
 FILLCELL_X4 FILLER_101_1143 ();
 FILLCELL_X1 FILLER_101_1147 ();
 FILLCELL_X1 FILLER_102_1 ();
 FILLCELL_X2 FILLER_102_26 ();
 FILLCELL_X1 FILLER_102_42 ();
 FILLCELL_X1 FILLER_102_75 ();
 FILLCELL_X4 FILLER_102_94 ();
 FILLCELL_X1 FILLER_102_98 ();
 FILLCELL_X16 FILLER_102_139 ();
 FILLCELL_X1 FILLER_102_155 ();
 FILLCELL_X4 FILLER_102_160 ();
 FILLCELL_X2 FILLER_102_182 ();
 FILLCELL_X1 FILLER_102_188 ();
 FILLCELL_X1 FILLER_102_313 ();
 FILLCELL_X2 FILLER_102_390 ();
 FILLCELL_X2 FILLER_102_429 ();
 FILLCELL_X1 FILLER_102_431 ();
 FILLCELL_X1 FILLER_102_436 ();
 FILLCELL_X1 FILLER_102_441 ();
 FILLCELL_X1 FILLER_102_452 ();
 FILLCELL_X2 FILLER_102_455 ();
 FILLCELL_X1 FILLER_102_474 ();
 FILLCELL_X2 FILLER_102_499 ();
 FILLCELL_X1 FILLER_102_567 ();
 FILLCELL_X1 FILLER_102_587 ();
 FILLCELL_X2 FILLER_102_616 ();
 FILLCELL_X1 FILLER_102_622 ();
 FILLCELL_X1 FILLER_102_630 ();
 FILLCELL_X2 FILLER_102_646 ();
 FILLCELL_X1 FILLER_102_648 ();
 FILLCELL_X2 FILLER_102_671 ();
 FILLCELL_X1 FILLER_102_673 ();
 FILLCELL_X1 FILLER_102_761 ();
 FILLCELL_X1 FILLER_102_912 ();
 FILLCELL_X1 FILLER_102_1020 ();
 FILLCELL_X2 FILLER_102_1036 ();
 FILLCELL_X1 FILLER_102_1090 ();
 FILLCELL_X16 FILLER_102_1132 ();
 FILLCELL_X2 FILLER_103_1 ();
 FILLCELL_X1 FILLER_103_3 ();
 FILLCELL_X1 FILLER_103_7 ();
 FILLCELL_X2 FILLER_103_30 ();
 FILLCELL_X2 FILLER_103_52 ();
 FILLCELL_X4 FILLER_103_70 ();
 FILLCELL_X2 FILLER_103_74 ();
 FILLCELL_X1 FILLER_103_76 ();
 FILLCELL_X2 FILLER_103_81 ();
 FILLCELL_X1 FILLER_103_83 ();
 FILLCELL_X2 FILLER_103_102 ();
 FILLCELL_X1 FILLER_103_104 ();
 FILLCELL_X8 FILLER_103_107 ();
 FILLCELL_X2 FILLER_103_115 ();
 FILLCELL_X8 FILLER_103_121 ();
 FILLCELL_X2 FILLER_103_129 ();
 FILLCELL_X1 FILLER_103_176 ();
 FILLCELL_X1 FILLER_103_187 ();
 FILLCELL_X1 FILLER_103_213 ();
 FILLCELL_X4 FILLER_103_234 ();
 FILLCELL_X2 FILLER_103_238 ();
 FILLCELL_X1 FILLER_103_240 ();
 FILLCELL_X2 FILLER_103_244 ();
 FILLCELL_X1 FILLER_103_246 ();
 FILLCELL_X4 FILLER_103_250 ();
 FILLCELL_X1 FILLER_103_254 ();
 FILLCELL_X2 FILLER_103_360 ();
 FILLCELL_X1 FILLER_103_447 ();
 FILLCELL_X1 FILLER_103_452 ();
 FILLCELL_X1 FILLER_103_457 ();
 FILLCELL_X1 FILLER_103_470 ();
 FILLCELL_X1 FILLER_103_474 ();
 FILLCELL_X1 FILLER_103_480 ();
 FILLCELL_X1 FILLER_103_485 ();
 FILLCELL_X1 FILLER_103_508 ();
 FILLCELL_X4 FILLER_103_532 ();
 FILLCELL_X2 FILLER_103_536 ();
 FILLCELL_X1 FILLER_103_538 ();
 FILLCELL_X4 FILLER_103_548 ();
 FILLCELL_X1 FILLER_103_585 ();
 FILLCELL_X2 FILLER_103_609 ();
 FILLCELL_X2 FILLER_103_622 ();
 FILLCELL_X8 FILLER_103_649 ();
 FILLCELL_X8 FILLER_103_660 ();
 FILLCELL_X4 FILLER_103_668 ();
 FILLCELL_X1 FILLER_103_686 ();
 FILLCELL_X1 FILLER_103_690 ();
 FILLCELL_X1 FILLER_103_697 ();
 FILLCELL_X1 FILLER_103_702 ();
 FILLCELL_X2 FILLER_103_707 ();
 FILLCELL_X1 FILLER_103_777 ();
 FILLCELL_X1 FILLER_103_785 ();
 FILLCELL_X8 FILLER_103_829 ();
 FILLCELL_X1 FILLER_103_837 ();
 FILLCELL_X1 FILLER_103_847 ();
 FILLCELL_X2 FILLER_103_860 ();
 FILLCELL_X2 FILLER_103_869 ();
 FILLCELL_X2 FILLER_103_923 ();
 FILLCELL_X1 FILLER_103_928 ();
 FILLCELL_X1 FILLER_103_951 ();
 FILLCELL_X2 FILLER_103_954 ();
 FILLCELL_X1 FILLER_103_956 ();
 FILLCELL_X4 FILLER_103_983 ();
 FILLCELL_X1 FILLER_103_1041 ();
 FILLCELL_X2 FILLER_103_1128 ();
 FILLCELL_X2 FILLER_103_1134 ();
 FILLCELL_X8 FILLER_103_1139 ();
 FILLCELL_X1 FILLER_103_1147 ();
 FILLCELL_X4 FILLER_104_1 ();
 FILLCELL_X2 FILLER_104_8 ();
 FILLCELL_X1 FILLER_104_14 ();
 FILLCELL_X2 FILLER_104_24 ();
 FILLCELL_X1 FILLER_104_26 ();
 FILLCELL_X1 FILLER_104_31 ();
 FILLCELL_X2 FILLER_104_42 ();
 FILLCELL_X1 FILLER_104_44 ();
 FILLCELL_X4 FILLER_104_47 ();
 FILLCELL_X1 FILLER_104_51 ();
 FILLCELL_X1 FILLER_104_54 ();
 FILLCELL_X4 FILLER_104_71 ();
 FILLCELL_X2 FILLER_104_75 ();
 FILLCELL_X1 FILLER_104_77 ();
 FILLCELL_X1 FILLER_104_85 ();
 FILLCELL_X1 FILLER_104_102 ();
 FILLCELL_X1 FILLER_104_119 ();
 FILLCELL_X1 FILLER_104_123 ();
 FILLCELL_X4 FILLER_104_127 ();
 FILLCELL_X1 FILLER_104_131 ();
 FILLCELL_X2 FILLER_104_136 ();
 FILLCELL_X4 FILLER_104_140 ();
 FILLCELL_X1 FILLER_104_144 ();
 FILLCELL_X2 FILLER_104_189 ();
 FILLCELL_X1 FILLER_104_221 ();
 FILLCELL_X2 FILLER_104_232 ();
 FILLCELL_X1 FILLER_104_234 ();
 FILLCELL_X4 FILLER_104_249 ();
 FILLCELL_X1 FILLER_104_253 ();
 FILLCELL_X1 FILLER_104_320 ();
 FILLCELL_X1 FILLER_104_354 ();
 FILLCELL_X1 FILLER_104_358 ();
 FILLCELL_X1 FILLER_104_366 ();
 FILLCELL_X1 FILLER_104_455 ();
 FILLCELL_X1 FILLER_104_536 ();
 FILLCELL_X4 FILLER_104_546 ();
 FILLCELL_X1 FILLER_104_550 ();
 FILLCELL_X4 FILLER_104_564 ();
 FILLCELL_X2 FILLER_104_568 ();
 FILLCELL_X1 FILLER_104_570 ();
 FILLCELL_X2 FILLER_104_603 ();
 FILLCELL_X1 FILLER_104_605 ();
 FILLCELL_X1 FILLER_104_613 ();
 FILLCELL_X2 FILLER_104_628 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X2 FILLER_104_638 ();
 FILLCELL_X1 FILLER_104_644 ();
 FILLCELL_X1 FILLER_104_648 ();
 FILLCELL_X2 FILLER_104_671 ();
 FILLCELL_X2 FILLER_104_692 ();
 FILLCELL_X1 FILLER_104_700 ();
 FILLCELL_X2 FILLER_104_707 ();
 FILLCELL_X2 FILLER_104_713 ();
 FILLCELL_X1 FILLER_104_788 ();
 FILLCELL_X1 FILLER_104_798 ();
 FILLCELL_X1 FILLER_104_806 ();
 FILLCELL_X2 FILLER_104_899 ();
 FILLCELL_X2 FILLER_104_934 ();
 FILLCELL_X2 FILLER_104_948 ();
 FILLCELL_X1 FILLER_104_1005 ();
 FILLCELL_X8 FILLER_104_1023 ();
 FILLCELL_X1 FILLER_104_1031 ();
 FILLCELL_X1 FILLER_104_1036 ();
 FILLCELL_X1 FILLER_104_1098 ();
 FILLCELL_X1 FILLER_104_1133 ();
 FILLCELL_X4 FILLER_104_1139 ();
 FILLCELL_X2 FILLER_104_1143 ();
 FILLCELL_X1 FILLER_105_9 ();
 FILLCELL_X1 FILLER_105_46 ();
 FILLCELL_X1 FILLER_105_63 ();
 FILLCELL_X1 FILLER_105_80 ();
 FILLCELL_X1 FILLER_105_97 ();
 FILLCELL_X1 FILLER_105_130 ();
 FILLCELL_X8 FILLER_105_151 ();
 FILLCELL_X4 FILLER_105_159 ();
 FILLCELL_X2 FILLER_105_183 ();
 FILLCELL_X1 FILLER_105_253 ();
 FILLCELL_X2 FILLER_105_328 ();
 FILLCELL_X1 FILLER_105_344 ();
 FILLCELL_X1 FILLER_105_348 ();
 FILLCELL_X2 FILLER_105_419 ();
 FILLCELL_X2 FILLER_105_472 ();
 FILLCELL_X1 FILLER_105_493 ();
 FILLCELL_X1 FILLER_105_501 ();
 FILLCELL_X1 FILLER_105_528 ();
 FILLCELL_X1 FILLER_105_562 ();
 FILLCELL_X8 FILLER_105_567 ();
 FILLCELL_X2 FILLER_105_575 ();
 FILLCELL_X2 FILLER_105_606 ();
 FILLCELL_X1 FILLER_105_608 ();
 FILLCELL_X1 FILLER_105_644 ();
 FILLCELL_X16 FILLER_105_651 ();
 FILLCELL_X4 FILLER_105_667 ();
 FILLCELL_X2 FILLER_105_671 ();
 FILLCELL_X1 FILLER_105_673 ();
 FILLCELL_X8 FILLER_105_681 ();
 FILLCELL_X1 FILLER_105_704 ();
 FILLCELL_X2 FILLER_105_774 ();
 FILLCELL_X1 FILLER_105_803 ();
 FILLCELL_X2 FILLER_105_874 ();
 FILLCELL_X1 FILLER_105_883 ();
 FILLCELL_X1 FILLER_105_890 ();
 FILLCELL_X2 FILLER_105_898 ();
 FILLCELL_X1 FILLER_105_932 ();
 FILLCELL_X2 FILLER_105_940 ();
 FILLCELL_X1 FILLER_105_949 ();
 FILLCELL_X1 FILLER_105_952 ();
 FILLCELL_X1 FILLER_105_963 ();
 FILLCELL_X1 FILLER_105_968 ();
 FILLCELL_X1 FILLER_105_975 ();
 FILLCELL_X1 FILLER_105_986 ();
 FILLCELL_X2 FILLER_105_996 ();
 FILLCELL_X1 FILLER_105_1053 ();
 FILLCELL_X8 FILLER_105_1058 ();
 FILLCELL_X1 FILLER_105_1066 ();
 FILLCELL_X4 FILLER_105_1133 ();
 FILLCELL_X2 FILLER_105_1137 ();
 FILLCELL_X4 FILLER_105_1142 ();
 FILLCELL_X2 FILLER_105_1146 ();
 FILLCELL_X2 FILLER_106_4 ();
 FILLCELL_X1 FILLER_106_6 ();
 FILLCELL_X1 FILLER_106_22 ();
 FILLCELL_X2 FILLER_106_43 ();
 FILLCELL_X1 FILLER_106_45 ();
 FILLCELL_X4 FILLER_106_48 ();
 FILLCELL_X1 FILLER_106_56 ();
 FILLCELL_X1 FILLER_106_59 ();
 FILLCELL_X1 FILLER_106_76 ();
 FILLCELL_X1 FILLER_106_79 ();
 FILLCELL_X2 FILLER_106_82 ();
 FILLCELL_X1 FILLER_106_84 ();
 FILLCELL_X2 FILLER_106_89 ();
 FILLCELL_X1 FILLER_106_91 ();
 FILLCELL_X1 FILLER_106_114 ();
 FILLCELL_X1 FILLER_106_131 ();
 FILLCELL_X2 FILLER_106_135 ();
 FILLCELL_X1 FILLER_106_163 ();
 FILLCELL_X4 FILLER_106_166 ();
 FILLCELL_X8 FILLER_106_174 ();
 FILLCELL_X4 FILLER_106_182 ();
 FILLCELL_X2 FILLER_106_186 ();
 FILLCELL_X1 FILLER_106_188 ();
 FILLCELL_X4 FILLER_106_193 ();
 FILLCELL_X2 FILLER_106_197 ();
 FILLCELL_X16 FILLER_106_209 ();
 FILLCELL_X4 FILLER_106_225 ();
 FILLCELL_X2 FILLER_106_236 ();
 FILLCELL_X1 FILLER_106_238 ();
 FILLCELL_X1 FILLER_106_242 ();
 FILLCELL_X2 FILLER_106_247 ();
 FILLCELL_X1 FILLER_106_252 ();
 FILLCELL_X2 FILLER_106_275 ();
 FILLCELL_X1 FILLER_106_314 ();
 FILLCELL_X1 FILLER_106_320 ();
 FILLCELL_X1 FILLER_106_413 ();
 FILLCELL_X1 FILLER_106_419 ();
 FILLCELL_X1 FILLER_106_429 ();
 FILLCELL_X1 FILLER_106_446 ();
 FILLCELL_X2 FILLER_106_455 ();
 FILLCELL_X1 FILLER_106_552 ();
 FILLCELL_X1 FILLER_106_560 ();
 FILLCELL_X2 FILLER_106_576 ();
 FILLCELL_X1 FILLER_106_578 ();
 FILLCELL_X2 FILLER_106_586 ();
 FILLCELL_X1 FILLER_106_588 ();
 FILLCELL_X8 FILLER_106_608 ();
 FILLCELL_X2 FILLER_106_616 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X2 FILLER_106_689 ();
 FILLCELL_X1 FILLER_106_691 ();
 FILLCELL_X2 FILLER_106_695 ();
 FILLCELL_X1 FILLER_106_697 ();
 FILLCELL_X1 FILLER_106_774 ();
 FILLCELL_X2 FILLER_106_820 ();
 FILLCELL_X2 FILLER_106_836 ();
 FILLCELL_X1 FILLER_106_865 ();
 FILLCELL_X1 FILLER_106_886 ();
 FILLCELL_X1 FILLER_106_894 ();
 FILLCELL_X1 FILLER_106_902 ();
 FILLCELL_X2 FILLER_106_917 ();
 FILLCELL_X1 FILLER_106_928 ();
 FILLCELL_X2 FILLER_106_961 ();
 FILLCELL_X2 FILLER_106_974 ();
 FILLCELL_X1 FILLER_106_976 ();
 FILLCELL_X1 FILLER_106_979 ();
 FILLCELL_X2 FILLER_106_1024 ();
 FILLCELL_X1 FILLER_106_1127 ();
 FILLCELL_X1 FILLER_107_5 ();
 FILLCELL_X4 FILLER_107_22 ();
 FILLCELL_X2 FILLER_107_26 ();
 FILLCELL_X4 FILLER_107_36 ();
 FILLCELL_X2 FILLER_107_40 ();
 FILLCELL_X1 FILLER_107_42 ();
 FILLCELL_X1 FILLER_107_51 ();
 FILLCELL_X4 FILLER_107_58 ();
 FILLCELL_X2 FILLER_107_62 ();
 FILLCELL_X1 FILLER_107_100 ();
 FILLCELL_X1 FILLER_107_109 ();
 FILLCELL_X4 FILLER_107_114 ();
 FILLCELL_X2 FILLER_107_118 ();
 FILLCELL_X1 FILLER_107_120 ();
 FILLCELL_X1 FILLER_107_157 ();
 FILLCELL_X1 FILLER_107_182 ();
 FILLCELL_X2 FILLER_107_203 ();
 FILLCELL_X2 FILLER_107_225 ();
 FILLCELL_X2 FILLER_107_236 ();
 FILLCELL_X1 FILLER_107_241 ();
 FILLCELL_X4 FILLER_107_246 ();
 FILLCELL_X2 FILLER_107_250 ();
 FILLCELL_X2 FILLER_107_276 ();
 FILLCELL_X1 FILLER_107_430 ();
 FILLCELL_X1 FILLER_107_460 ();
 FILLCELL_X1 FILLER_107_501 ();
 FILLCELL_X1 FILLER_107_507 ();
 FILLCELL_X1 FILLER_107_524 ();
 FILLCELL_X4 FILLER_107_593 ();
 FILLCELL_X1 FILLER_107_607 ();
 FILLCELL_X4 FILLER_107_618 ();
 FILLCELL_X1 FILLER_107_631 ();
 FILLCELL_X8 FILLER_107_660 ();
 FILLCELL_X1 FILLER_107_668 ();
 FILLCELL_X8 FILLER_107_718 ();
 FILLCELL_X4 FILLER_107_726 ();
 FILLCELL_X2 FILLER_107_730 ();
 FILLCELL_X1 FILLER_107_736 ();
 FILLCELL_X4 FILLER_107_785 ();
 FILLCELL_X1 FILLER_107_789 ();
 FILLCELL_X1 FILLER_107_847 ();
 FILLCELL_X1 FILLER_107_861 ();
 FILLCELL_X1 FILLER_107_885 ();
 FILLCELL_X1 FILLER_107_896 ();
 FILLCELL_X1 FILLER_107_904 ();
 FILLCELL_X1 FILLER_107_912 ();
 FILLCELL_X2 FILLER_107_928 ();
 FILLCELL_X1 FILLER_107_930 ();
 FILLCELL_X1 FILLER_107_938 ();
 FILLCELL_X1 FILLER_107_985 ();
 FILLCELL_X1 FILLER_107_1030 ();
 FILLCELL_X1 FILLER_107_1059 ();
 FILLCELL_X1 FILLER_107_1112 ();
 FILLCELL_X4 FILLER_107_1137 ();
 FILLCELL_X1 FILLER_107_1141 ();
 FILLCELL_X2 FILLER_108_1 ();
 FILLCELL_X1 FILLER_108_3 ();
 FILLCELL_X2 FILLER_108_20 ();
 FILLCELL_X1 FILLER_108_24 ();
 FILLCELL_X1 FILLER_108_28 ();
 FILLCELL_X1 FILLER_108_32 ();
 FILLCELL_X1 FILLER_108_40 ();
 FILLCELL_X1 FILLER_108_57 ();
 FILLCELL_X2 FILLER_108_79 ();
 FILLCELL_X1 FILLER_108_84 ();
 FILLCELL_X2 FILLER_108_89 ();
 FILLCELL_X1 FILLER_108_95 ();
 FILLCELL_X1 FILLER_108_112 ();
 FILLCELL_X2 FILLER_108_115 ();
 FILLCELL_X2 FILLER_108_206 ();
 FILLCELL_X2 FILLER_108_251 ();
 FILLCELL_X8 FILLER_108_257 ();
 FILLCELL_X4 FILLER_108_265 ();
 FILLCELL_X2 FILLER_108_269 ();
 FILLCELL_X1 FILLER_108_271 ();
 FILLCELL_X1 FILLER_108_340 ();
 FILLCELL_X1 FILLER_108_380 ();
 FILLCELL_X2 FILLER_108_424 ();
 FILLCELL_X1 FILLER_108_428 ();
 FILLCELL_X1 FILLER_108_486 ();
 FILLCELL_X1 FILLER_108_491 ();
 FILLCELL_X2 FILLER_108_507 ();
 FILLCELL_X2 FILLER_108_600 ();
 FILLCELL_X2 FILLER_108_619 ();
 FILLCELL_X1 FILLER_108_621 ();
 FILLCELL_X1 FILLER_108_630 ();
 FILLCELL_X1 FILLER_108_647 ();
 FILLCELL_X1 FILLER_108_654 ();
 FILLCELL_X1 FILLER_108_675 ();
 FILLCELL_X1 FILLER_108_679 ();
 FILLCELL_X1 FILLER_108_686 ();
 FILLCELL_X1 FILLER_108_692 ();
 FILLCELL_X1 FILLER_108_804 ();
 FILLCELL_X1 FILLER_108_818 ();
 FILLCELL_X1 FILLER_108_870 ();
 FILLCELL_X2 FILLER_108_874 ();
 FILLCELL_X4 FILLER_108_883 ();
 FILLCELL_X2 FILLER_108_901 ();
 FILLCELL_X1 FILLER_108_903 ();
 FILLCELL_X2 FILLER_108_913 ();
 FILLCELL_X1 FILLER_108_915 ();
 FILLCELL_X1 FILLER_108_931 ();
 FILLCELL_X2 FILLER_108_1038 ();
 FILLCELL_X1 FILLER_108_1046 ();
 FILLCELL_X2 FILLER_108_1063 ();
 FILLCELL_X2 FILLER_108_1079 ();
 FILLCELL_X2 FILLER_108_1090 ();
 FILLCELL_X2 FILLER_108_1126 ();
 FILLCELL_X1 FILLER_109_9 ();
 FILLCELL_X1 FILLER_109_32 ();
 FILLCELL_X4 FILLER_109_36 ();
 FILLCELL_X4 FILLER_109_43 ();
 FILLCELL_X2 FILLER_109_59 ();
 FILLCELL_X1 FILLER_109_61 ();
 FILLCELL_X2 FILLER_109_70 ();
 FILLCELL_X1 FILLER_109_72 ();
 FILLCELL_X2 FILLER_109_76 ();
 FILLCELL_X2 FILLER_109_82 ();
 FILLCELL_X1 FILLER_109_94 ();
 FILLCELL_X4 FILLER_109_105 ();
 FILLCELL_X1 FILLER_109_109 ();
 FILLCELL_X8 FILLER_109_176 ();
 FILLCELL_X8 FILLER_109_209 ();
 FILLCELL_X2 FILLER_109_217 ();
 FILLCELL_X1 FILLER_109_219 ();
 FILLCELL_X1 FILLER_109_226 ();
 FILLCELL_X1 FILLER_109_273 ();
 FILLCELL_X1 FILLER_109_379 ();
 FILLCELL_X1 FILLER_109_384 ();
 FILLCELL_X2 FILLER_109_405 ();
 FILLCELL_X1 FILLER_109_432 ();
 FILLCELL_X1 FILLER_109_502 ();
 FILLCELL_X1 FILLER_109_528 ();
 FILLCELL_X1 FILLER_109_537 ();
 FILLCELL_X2 FILLER_109_566 ();
 FILLCELL_X1 FILLER_109_568 ();
 FILLCELL_X2 FILLER_109_576 ();
 FILLCELL_X2 FILLER_109_652 ();
 FILLCELL_X1 FILLER_109_654 ();
 FILLCELL_X4 FILLER_109_681 ();
 FILLCELL_X2 FILLER_109_694 ();
 FILLCELL_X1 FILLER_109_746 ();
 FILLCELL_X1 FILLER_109_752 ();
 FILLCELL_X1 FILLER_109_764 ();
 FILLCELL_X1 FILLER_109_785 ();
 FILLCELL_X1 FILLER_109_797 ();
 FILLCELL_X1 FILLER_109_845 ();
 FILLCELL_X1 FILLER_109_941 ();
 FILLCELL_X1 FILLER_109_993 ();
 FILLCELL_X1 FILLER_109_1028 ();
 FILLCELL_X1 FILLER_109_1069 ();
 FILLCELL_X1 FILLER_109_1075 ();
 FILLCELL_X1 FILLER_109_1092 ();
 FILLCELL_X2 FILLER_109_1102 ();
 FILLCELL_X1 FILLER_109_1104 ();
 FILLCELL_X2 FILLER_109_1116 ();
 FILLCELL_X8 FILLER_109_1136 ();
 FILLCELL_X1 FILLER_109_1144 ();
 FILLCELL_X2 FILLER_110_1 ();
 FILLCELL_X1 FILLER_110_3 ();
 FILLCELL_X2 FILLER_110_39 ();
 FILLCELL_X8 FILLER_110_43 ();
 FILLCELL_X1 FILLER_110_51 ();
 FILLCELL_X1 FILLER_110_57 ();
 FILLCELL_X1 FILLER_110_66 ();
 FILLCELL_X4 FILLER_110_86 ();
 FILLCELL_X2 FILLER_110_93 ();
 FILLCELL_X1 FILLER_110_99 ();
 FILLCELL_X1 FILLER_110_118 ();
 FILLCELL_X4 FILLER_110_123 ();
 FILLCELL_X2 FILLER_110_127 ();
 FILLCELL_X4 FILLER_110_131 ();
 FILLCELL_X1 FILLER_110_135 ();
 FILLCELL_X4 FILLER_110_140 ();
 FILLCELL_X16 FILLER_110_188 ();
 FILLCELL_X4 FILLER_110_204 ();
 FILLCELL_X2 FILLER_110_409 ();
 FILLCELL_X2 FILLER_110_592 ();
 FILLCELL_X1 FILLER_110_615 ();
 FILLCELL_X1 FILLER_110_630 ();
 FILLCELL_X1 FILLER_110_646 ();
 FILLCELL_X1 FILLER_110_650 ();
 FILLCELL_X8 FILLER_110_659 ();
 FILLCELL_X4 FILLER_110_667 ();
 FILLCELL_X1 FILLER_110_679 ();
 FILLCELL_X2 FILLER_110_683 ();
 FILLCELL_X1 FILLER_110_685 ();
 FILLCELL_X8 FILLER_110_705 ();
 FILLCELL_X2 FILLER_110_713 ();
 FILLCELL_X4 FILLER_110_737 ();
 FILLCELL_X2 FILLER_110_741 ();
 FILLCELL_X1 FILLER_110_852 ();
 FILLCELL_X2 FILLER_110_866 ();
 FILLCELL_X1 FILLER_110_868 ();
 FILLCELL_X8 FILLER_110_875 ();
 FILLCELL_X1 FILLER_110_883 ();
 FILLCELL_X2 FILLER_110_897 ();
 FILLCELL_X2 FILLER_110_931 ();
 FILLCELL_X1 FILLER_110_933 ();
 FILLCELL_X2 FILLER_110_943 ();
 FILLCELL_X1 FILLER_110_945 ();
 FILLCELL_X1 FILLER_110_950 ();
 FILLCELL_X2 FILLER_110_1018 ();
 FILLCELL_X1 FILLER_110_1040 ();
 FILLCELL_X8 FILLER_110_1137 ();
 FILLCELL_X2 FILLER_110_1145 ();
 FILLCELL_X1 FILLER_110_1147 ();
 FILLCELL_X1 FILLER_111_14 ();
 FILLCELL_X2 FILLER_111_37 ();
 FILLCELL_X1 FILLER_111_59 ();
 FILLCELL_X1 FILLER_111_62 ();
 FILLCELL_X1 FILLER_111_66 ();
 FILLCELL_X1 FILLER_111_71 ();
 FILLCELL_X1 FILLER_111_126 ();
 FILLCELL_X8 FILLER_111_167 ();
 FILLCELL_X2 FILLER_111_175 ();
 FILLCELL_X8 FILLER_111_187 ();
 FILLCELL_X2 FILLER_111_195 ();
 FILLCELL_X1 FILLER_111_197 ();
 FILLCELL_X1 FILLER_111_212 ();
 FILLCELL_X8 FILLER_111_217 ();
 FILLCELL_X1 FILLER_111_225 ();
 FILLCELL_X4 FILLER_111_236 ();
 FILLCELL_X2 FILLER_111_253 ();
 FILLCELL_X2 FILLER_111_257 ();
 FILLCELL_X4 FILLER_111_332 ();
 FILLCELL_X1 FILLER_111_357 ();
 FILLCELL_X2 FILLER_111_361 ();
 FILLCELL_X1 FILLER_111_363 ();
 FILLCELL_X2 FILLER_111_445 ();
 FILLCELL_X1 FILLER_111_492 ();
 FILLCELL_X2 FILLER_111_519 ();
 FILLCELL_X1 FILLER_111_607 ();
 FILLCELL_X2 FILLER_111_613 ();
 FILLCELL_X2 FILLER_111_640 ();
 FILLCELL_X1 FILLER_111_642 ();
 FILLCELL_X2 FILLER_111_730 ();
 FILLCELL_X2 FILLER_111_797 ();
 FILLCELL_X1 FILLER_111_799 ();
 FILLCELL_X1 FILLER_111_810 ();
 FILLCELL_X1 FILLER_111_826 ();
 FILLCELL_X1 FILLER_111_873 ();
 FILLCELL_X2 FILLER_111_877 ();
 FILLCELL_X1 FILLER_111_894 ();
 FILLCELL_X2 FILLER_111_908 ();
 FILLCELL_X1 FILLER_111_910 ();
 FILLCELL_X2 FILLER_111_964 ();
 FILLCELL_X2 FILLER_111_1014 ();
 FILLCELL_X1 FILLER_111_1058 ();
 FILLCELL_X2 FILLER_111_1091 ();
 FILLCELL_X4 FILLER_111_1124 ();
 FILLCELL_X16 FILLER_111_1131 ();
 FILLCELL_X1 FILLER_111_1147 ();
 FILLCELL_X1 FILLER_112_49 ();
 FILLCELL_X1 FILLER_112_54 ();
 FILLCELL_X2 FILLER_112_75 ();
 FILLCELL_X1 FILLER_112_77 ();
 FILLCELL_X1 FILLER_112_81 ();
 FILLCELL_X4 FILLER_112_88 ();
 FILLCELL_X2 FILLER_112_92 ();
 FILLCELL_X4 FILLER_112_110 ();
 FILLCELL_X2 FILLER_112_114 ();
 FILLCELL_X2 FILLER_112_119 ();
 FILLCELL_X1 FILLER_112_121 ();
 FILLCELL_X2 FILLER_112_128 ();
 FILLCELL_X4 FILLER_112_134 ();
 FILLCELL_X8 FILLER_112_158 ();
 FILLCELL_X4 FILLER_112_166 ();
 FILLCELL_X2 FILLER_112_170 ();
 FILLCELL_X8 FILLER_112_182 ();
 FILLCELL_X4 FILLER_112_194 ();
 FILLCELL_X1 FILLER_112_198 ();
 FILLCELL_X2 FILLER_112_207 ();
 FILLCELL_X1 FILLER_112_233 ();
 FILLCELL_X4 FILLER_112_238 ();
 FILLCELL_X1 FILLER_112_244 ();
 FILLCELL_X1 FILLER_112_251 ();
 FILLCELL_X1 FILLER_112_351 ();
 FILLCELL_X1 FILLER_112_392 ();
 FILLCELL_X1 FILLER_112_432 ();
 FILLCELL_X1 FILLER_112_455 ();
 FILLCELL_X1 FILLER_112_538 ();
 FILLCELL_X2 FILLER_112_560 ();
 FILLCELL_X1 FILLER_112_614 ();
 FILLCELL_X2 FILLER_112_628 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X2 FILLER_112_635 ();
 FILLCELL_X1 FILLER_112_637 ();
 FILLCELL_X2 FILLER_112_681 ();
 FILLCELL_X8 FILLER_112_689 ();
 FILLCELL_X2 FILLER_112_697 ();
 FILLCELL_X1 FILLER_112_702 ();
 FILLCELL_X1 FILLER_112_708 ();
 FILLCELL_X2 FILLER_112_712 ();
 FILLCELL_X2 FILLER_112_734 ();
 FILLCELL_X1 FILLER_112_740 ();
 FILLCELL_X4 FILLER_112_749 ();
 FILLCELL_X2 FILLER_112_753 ();
 FILLCELL_X1 FILLER_112_755 ();
 FILLCELL_X2 FILLER_112_786 ();
 FILLCELL_X1 FILLER_112_788 ();
 FILLCELL_X2 FILLER_112_809 ();
 FILLCELL_X1 FILLER_112_821 ();
 FILLCELL_X1 FILLER_112_864 ();
 FILLCELL_X4 FILLER_112_868 ();
 FILLCELL_X1 FILLER_112_876 ();
 FILLCELL_X2 FILLER_112_893 ();
 FILLCELL_X1 FILLER_112_895 ();
 FILLCELL_X4 FILLER_112_900 ();
 FILLCELL_X8 FILLER_112_909 ();
 FILLCELL_X4 FILLER_112_917 ();
 FILLCELL_X2 FILLER_112_979 ();
 FILLCELL_X2 FILLER_112_1011 ();
 FILLCELL_X1 FILLER_112_1026 ();
 FILLCELL_X1 FILLER_112_1053 ();
 FILLCELL_X2 FILLER_112_1067 ();
 FILLCELL_X1 FILLER_112_1075 ();
 FILLCELL_X4 FILLER_112_1108 ();
 FILLCELL_X8 FILLER_112_1134 ();
 FILLCELL_X4 FILLER_112_1142 ();
 FILLCELL_X2 FILLER_112_1146 ();
 FILLCELL_X1 FILLER_113_38 ();
 FILLCELL_X1 FILLER_113_41 ();
 FILLCELL_X1 FILLER_113_74 ();
 FILLCELL_X2 FILLER_113_78 ();
 FILLCELL_X1 FILLER_113_84 ();
 FILLCELL_X2 FILLER_113_89 ();
 FILLCELL_X4 FILLER_113_107 ();
 FILLCELL_X2 FILLER_113_111 ();
 FILLCELL_X1 FILLER_113_113 ();
 FILLCELL_X4 FILLER_113_121 ();
 FILLCELL_X2 FILLER_113_139 ();
 FILLCELL_X1 FILLER_113_144 ();
 FILLCELL_X4 FILLER_113_180 ();
 FILLCELL_X2 FILLER_113_184 ();
 FILLCELL_X4 FILLER_113_190 ();
 FILLCELL_X1 FILLER_113_220 ();
 FILLCELL_X1 FILLER_113_236 ();
 FILLCELL_X2 FILLER_113_243 ();
 FILLCELL_X2 FILLER_113_254 ();
 FILLCELL_X1 FILLER_113_256 ();
 FILLCELL_X2 FILLER_113_348 ();
 FILLCELL_X1 FILLER_113_368 ();
 FILLCELL_X2 FILLER_113_419 ();
 FILLCELL_X2 FILLER_113_430 ();
 FILLCELL_X1 FILLER_113_432 ();
 FILLCELL_X1 FILLER_113_550 ();
 FILLCELL_X1 FILLER_113_628 ();
 FILLCELL_X2 FILLER_113_668 ();
 FILLCELL_X2 FILLER_113_691 ();
 FILLCELL_X1 FILLER_113_693 ();
 FILLCELL_X4 FILLER_113_701 ();
 FILLCELL_X2 FILLER_113_705 ();
 FILLCELL_X2 FILLER_113_869 ();
 FILLCELL_X2 FILLER_113_874 ();
 FILLCELL_X1 FILLER_113_876 ();
 FILLCELL_X4 FILLER_113_883 ();
 FILLCELL_X2 FILLER_113_887 ();
 FILLCELL_X8 FILLER_113_901 ();
 FILLCELL_X4 FILLER_113_909 ();
 FILLCELL_X2 FILLER_113_913 ();
 FILLCELL_X1 FILLER_113_915 ();
 FILLCELL_X1 FILLER_113_1070 ();
 FILLCELL_X1 FILLER_113_1074 ();
 FILLCELL_X4 FILLER_113_1118 ();
 FILLCELL_X2 FILLER_113_1124 ();
 FILLCELL_X4 FILLER_113_1132 ();
 FILLCELL_X1 FILLER_113_1136 ();
 FILLCELL_X4 FILLER_113_1141 ();
 FILLCELL_X2 FILLER_113_1145 ();
 FILLCELL_X1 FILLER_113_1147 ();
 FILLCELL_X2 FILLER_114_22 ();
 FILLCELL_X1 FILLER_114_42 ();
 FILLCELL_X1 FILLER_114_45 ();
 FILLCELL_X1 FILLER_114_50 ();
 FILLCELL_X1 FILLER_114_55 ();
 FILLCELL_X2 FILLER_114_58 ();
 FILLCELL_X1 FILLER_114_60 ();
 FILLCELL_X4 FILLER_114_69 ();
 FILLCELL_X1 FILLER_114_73 ();
 FILLCELL_X4 FILLER_114_95 ();
 FILLCELL_X2 FILLER_114_99 ();
 FILLCELL_X1 FILLER_114_101 ();
 FILLCELL_X1 FILLER_114_104 ();
 FILLCELL_X2 FILLER_114_107 ();
 FILLCELL_X4 FILLER_114_174 ();
 FILLCELL_X1 FILLER_114_192 ();
 FILLCELL_X1 FILLER_114_205 ();
 FILLCELL_X2 FILLER_114_242 ();
 FILLCELL_X1 FILLER_114_268 ();
 FILLCELL_X4 FILLER_114_434 ();
 FILLCELL_X4 FILLER_114_462 ();
 FILLCELL_X1 FILLER_114_466 ();
 FILLCELL_X1 FILLER_114_503 ();
 FILLCELL_X1 FILLER_114_515 ();
 FILLCELL_X1 FILLER_114_520 ();
 FILLCELL_X1 FILLER_114_528 ();
 FILLCELL_X1 FILLER_114_541 ();
 FILLCELL_X1 FILLER_114_559 ();
 FILLCELL_X4 FILLER_114_632 ();
 FILLCELL_X2 FILLER_114_636 ();
 FILLCELL_X1 FILLER_114_640 ();
 FILLCELL_X1 FILLER_114_651 ();
 FILLCELL_X4 FILLER_114_674 ();
 FILLCELL_X8 FILLER_114_685 ();
 FILLCELL_X2 FILLER_114_693 ();
 FILLCELL_X1 FILLER_114_695 ();
 FILLCELL_X8 FILLER_114_712 ();
 FILLCELL_X2 FILLER_114_720 ();
 FILLCELL_X1 FILLER_114_722 ();
 FILLCELL_X1 FILLER_114_814 ();
 FILLCELL_X2 FILLER_114_821 ();
 FILLCELL_X4 FILLER_114_829 ();
 FILLCELL_X2 FILLER_114_833 ();
 FILLCELL_X8 FILLER_114_855 ();
 FILLCELL_X2 FILLER_114_863 ();
 FILLCELL_X1 FILLER_114_865 ();
 FILLCELL_X16 FILLER_114_869 ();
 FILLCELL_X4 FILLER_114_885 ();
 FILLCELL_X1 FILLER_114_889 ();
 FILLCELL_X4 FILLER_114_910 ();
 FILLCELL_X1 FILLER_114_914 ();
 FILLCELL_X1 FILLER_114_993 ();
 FILLCELL_X2 FILLER_114_1013 ();
 FILLCELL_X2 FILLER_114_1021 ();
 FILLCELL_X2 FILLER_114_1025 ();
 FILLCELL_X4 FILLER_114_1050 ();
 FILLCELL_X2 FILLER_114_1054 ();
 FILLCELL_X16 FILLER_114_1082 ();
 FILLCELL_X1 FILLER_114_1098 ();
 FILLCELL_X2 FILLER_114_1102 ();
 FILLCELL_X1 FILLER_114_1117 ();
 FILLCELL_X1 FILLER_114_1147 ();
 FILLCELL_X4 FILLER_115_4 ();
 FILLCELL_X2 FILLER_115_8 ();
 FILLCELL_X2 FILLER_115_18 ();
 FILLCELL_X1 FILLER_115_36 ();
 FILLCELL_X2 FILLER_115_53 ();
 FILLCELL_X1 FILLER_115_55 ();
 FILLCELL_X2 FILLER_115_72 ();
 FILLCELL_X1 FILLER_115_74 ();
 FILLCELL_X4 FILLER_115_93 ();
 FILLCELL_X1 FILLER_115_97 ();
 FILLCELL_X4 FILLER_115_106 ();
 FILLCELL_X1 FILLER_115_170 ();
 FILLCELL_X4 FILLER_115_181 ();
 FILLCELL_X2 FILLER_115_222 ();
 FILLCELL_X1 FILLER_115_230 ();
 FILLCELL_X1 FILLER_115_247 ();
 FILLCELL_X1 FILLER_115_253 ();
 FILLCELL_X2 FILLER_115_290 ();
 FILLCELL_X1 FILLER_115_303 ();
 FILLCELL_X2 FILLER_115_335 ();
 FILLCELL_X1 FILLER_115_367 ();
 FILLCELL_X1 FILLER_115_401 ();
 FILLCELL_X1 FILLER_115_500 ();
 FILLCELL_X1 FILLER_115_532 ();
 FILLCELL_X1 FILLER_115_543 ();
 FILLCELL_X1 FILLER_115_549 ();
 FILLCELL_X1 FILLER_115_581 ();
 FILLCELL_X1 FILLER_115_604 ();
 FILLCELL_X2 FILLER_115_613 ();
 FILLCELL_X8 FILLER_115_623 ();
 FILLCELL_X2 FILLER_115_631 ();
 FILLCELL_X1 FILLER_115_633 ();
 FILLCELL_X2 FILLER_115_675 ();
 FILLCELL_X4 FILLER_115_711 ();
 FILLCELL_X2 FILLER_115_715 ();
 FILLCELL_X1 FILLER_115_739 ();
 FILLCELL_X1 FILLER_115_742 ();
 FILLCELL_X1 FILLER_115_756 ();
 FILLCELL_X2 FILLER_115_767 ();
 FILLCELL_X1 FILLER_115_775 ();
 FILLCELL_X1 FILLER_115_778 ();
 FILLCELL_X1 FILLER_115_781 ();
 FILLCELL_X1 FILLER_115_784 ();
 FILLCELL_X1 FILLER_115_814 ();
 FILLCELL_X2 FILLER_115_835 ();
 FILLCELL_X1 FILLER_115_837 ();
 FILLCELL_X2 FILLER_115_856 ();
 FILLCELL_X1 FILLER_115_858 ();
 FILLCELL_X1 FILLER_115_862 ();
 FILLCELL_X2 FILLER_115_878 ();
 FILLCELL_X1 FILLER_115_880 ();
 FILLCELL_X1 FILLER_115_901 ();
 FILLCELL_X2 FILLER_115_924 ();
 FILLCELL_X2 FILLER_115_1011 ();
 FILLCELL_X1 FILLER_115_1067 ();
 FILLCELL_X1 FILLER_115_1074 ();
 FILLCELL_X1 FILLER_115_1086 ();
 FILLCELL_X2 FILLER_115_1105 ();
 FILLCELL_X2 FILLER_115_1112 ();
 FILLCELL_X1 FILLER_115_1114 ();
 FILLCELL_X2 FILLER_115_1118 ();
 FILLCELL_X1 FILLER_115_1120 ();
 FILLCELL_X1 FILLER_115_1124 ();
 FILLCELL_X1 FILLER_115_1129 ();
 FILLCELL_X2 FILLER_115_1135 ();
 FILLCELL_X1 FILLER_115_1141 ();
 FILLCELL_X2 FILLER_115_1146 ();
 FILLCELL_X4 FILLER_116_4 ();
 FILLCELL_X4 FILLER_116_18 ();
 FILLCELL_X1 FILLER_116_24 ();
 FILLCELL_X2 FILLER_116_41 ();
 FILLCELL_X4 FILLER_116_59 ();
 FILLCELL_X2 FILLER_116_63 ();
 FILLCELL_X1 FILLER_116_65 ();
 FILLCELL_X4 FILLER_116_114 ();
 FILLCELL_X2 FILLER_116_118 ();
 FILLCELL_X1 FILLER_116_120 ();
 FILLCELL_X4 FILLER_116_125 ();
 FILLCELL_X1 FILLER_116_196 ();
 FILLCELL_X2 FILLER_116_204 ();
 FILLCELL_X1 FILLER_116_309 ();
 FILLCELL_X1 FILLER_116_317 ();
 FILLCELL_X1 FILLER_116_337 ();
 FILLCELL_X2 FILLER_116_358 ();
 FILLCELL_X2 FILLER_116_430 ();
 FILLCELL_X1 FILLER_116_432 ();
 FILLCELL_X4 FILLER_116_525 ();
 FILLCELL_X2 FILLER_116_529 ();
 FILLCELL_X1 FILLER_116_534 ();
 FILLCELL_X1 FILLER_116_548 ();
 FILLCELL_X4 FILLER_116_632 ();
 FILLCELL_X1 FILLER_116_636 ();
 FILLCELL_X2 FILLER_116_644 ();
 FILLCELL_X1 FILLER_116_646 ();
 FILLCELL_X1 FILLER_116_671 ();
 FILLCELL_X2 FILLER_116_684 ();
 FILLCELL_X1 FILLER_116_686 ();
 FILLCELL_X2 FILLER_116_710 ();
 FILLCELL_X2 FILLER_116_752 ();
 FILLCELL_X2 FILLER_116_760 ();
 FILLCELL_X1 FILLER_116_762 ();
 FILLCELL_X2 FILLER_116_773 ();
 FILLCELL_X2 FILLER_116_803 ();
 FILLCELL_X1 FILLER_116_805 ();
 FILLCELL_X2 FILLER_116_816 ();
 FILLCELL_X2 FILLER_116_825 ();
 FILLCELL_X1 FILLER_116_827 ();
 FILLCELL_X2 FILLER_116_830 ();
 FILLCELL_X2 FILLER_116_838 ();
 FILLCELL_X1 FILLER_116_840 ();
 FILLCELL_X2 FILLER_116_847 ();
 FILLCELL_X1 FILLER_116_849 ();
 FILLCELL_X2 FILLER_116_854 ();
 FILLCELL_X1 FILLER_116_856 ();
 FILLCELL_X1 FILLER_116_864 ();
 FILLCELL_X2 FILLER_116_875 ();
 FILLCELL_X1 FILLER_116_877 ();
 FILLCELL_X1 FILLER_116_963 ();
 FILLCELL_X1 FILLER_116_973 ();
 FILLCELL_X2 FILLER_116_992 ();
 FILLCELL_X2 FILLER_116_1049 ();
 FILLCELL_X1 FILLER_116_1051 ();
 FILLCELL_X2 FILLER_116_1059 ();
 FILLCELL_X4 FILLER_116_1064 ();
 FILLCELL_X1 FILLER_116_1068 ();
 FILLCELL_X1 FILLER_116_1072 ();
 FILLCELL_X1 FILLER_116_1092 ();
 FILLCELL_X4 FILLER_116_1100 ();
 FILLCELL_X1 FILLER_116_1104 ();
 FILLCELL_X1 FILLER_116_1120 ();
 FILLCELL_X1 FILLER_116_1124 ();
 FILLCELL_X8 FILLER_116_1138 ();
 FILLCELL_X2 FILLER_116_1146 ();
 FILLCELL_X1 FILLER_117_27 ();
 FILLCELL_X1 FILLER_117_31 ();
 FILLCELL_X2 FILLER_117_52 ();
 FILLCELL_X2 FILLER_117_84 ();
 FILLCELL_X8 FILLER_117_102 ();
 FILLCELL_X4 FILLER_117_110 ();
 FILLCELL_X2 FILLER_117_114 ();
 FILLCELL_X1 FILLER_117_116 ();
 FILLCELL_X2 FILLER_117_119 ();
 FILLCELL_X8 FILLER_117_125 ();
 FILLCELL_X1 FILLER_117_133 ();
 FILLCELL_X2 FILLER_117_136 ();
 FILLCELL_X1 FILLER_117_138 ();
 FILLCELL_X4 FILLER_117_159 ();
 FILLCELL_X1 FILLER_117_163 ();
 FILLCELL_X8 FILLER_117_184 ();
 FILLCELL_X4 FILLER_117_192 ();
 FILLCELL_X1 FILLER_117_206 ();
 FILLCELL_X1 FILLER_117_211 ();
 FILLCELL_X4 FILLER_117_232 ();
 FILLCELL_X2 FILLER_117_239 ();
 FILLCELL_X2 FILLER_117_244 ();
 FILLCELL_X2 FILLER_117_264 ();
 FILLCELL_X1 FILLER_117_339 ();
 FILLCELL_X1 FILLER_117_354 ();
 FILLCELL_X4 FILLER_117_435 ();
 FILLCELL_X1 FILLER_117_446 ();
 FILLCELL_X2 FILLER_117_478 ();
 FILLCELL_X1 FILLER_117_542 ();
 FILLCELL_X2 FILLER_117_611 ();
 FILLCELL_X1 FILLER_117_643 ();
 FILLCELL_X2 FILLER_117_671 ();
 FILLCELL_X1 FILLER_117_673 ();
 FILLCELL_X2 FILLER_117_676 ();
 FILLCELL_X1 FILLER_117_682 ();
 FILLCELL_X2 FILLER_117_708 ();
 FILLCELL_X8 FILLER_117_712 ();
 FILLCELL_X4 FILLER_117_720 ();
 FILLCELL_X1 FILLER_117_724 ();
 FILLCELL_X4 FILLER_117_777 ();
 FILLCELL_X1 FILLER_117_849 ();
 FILLCELL_X1 FILLER_117_866 ();
 FILLCELL_X1 FILLER_117_920 ();
 FILLCELL_X1 FILLER_117_941 ();
 FILLCELL_X4 FILLER_117_1038 ();
 FILLCELL_X1 FILLER_117_1042 ();
 FILLCELL_X8 FILLER_117_1047 ();
 FILLCELL_X2 FILLER_117_1055 ();
 FILLCELL_X1 FILLER_117_1060 ();
 FILLCELL_X1 FILLER_117_1068 ();
 FILLCELL_X1 FILLER_117_1073 ();
 FILLCELL_X1 FILLER_117_1082 ();
 FILLCELL_X2 FILLER_117_1086 ();
 FILLCELL_X1 FILLER_117_1092 ();
 FILLCELL_X2 FILLER_117_1097 ();
 FILLCELL_X4 FILLER_117_1112 ();
 FILLCELL_X2 FILLER_117_1116 ();
 FILLCELL_X1 FILLER_117_1118 ();
 FILLCELL_X8 FILLER_117_1139 ();
 FILLCELL_X1 FILLER_117_1147 ();
 FILLCELL_X2 FILLER_118_18 ();
 FILLCELL_X2 FILLER_118_36 ();
 FILLCELL_X1 FILLER_118_38 ();
 FILLCELL_X1 FILLER_118_42 ();
 FILLCELL_X4 FILLER_118_45 ();
 FILLCELL_X2 FILLER_118_49 ();
 FILLCELL_X1 FILLER_118_51 ();
 FILLCELL_X2 FILLER_118_84 ();
 FILLCELL_X2 FILLER_118_88 ();
 FILLCELL_X1 FILLER_118_90 ();
 FILLCELL_X1 FILLER_118_107 ();
 FILLCELL_X1 FILLER_118_124 ();
 FILLCELL_X4 FILLER_118_135 ();
 FILLCELL_X2 FILLER_118_139 ();
 FILLCELL_X4 FILLER_118_143 ();
 FILLCELL_X2 FILLER_118_147 ();
 FILLCELL_X1 FILLER_118_149 ();
 FILLCELL_X4 FILLER_118_170 ();
 FILLCELL_X1 FILLER_118_194 ();
 FILLCELL_X1 FILLER_118_205 ();
 FILLCELL_X2 FILLER_118_242 ();
 FILLCELL_X1 FILLER_118_244 ();
 FILLCELL_X1 FILLER_118_251 ();
 FILLCELL_X2 FILLER_118_256 ();
 FILLCELL_X1 FILLER_118_258 ();
 FILLCELL_X1 FILLER_118_391 ();
 FILLCELL_X1 FILLER_118_519 ();
 FILLCELL_X1 FILLER_118_535 ();
 FILLCELL_X1 FILLER_118_547 ();
 FILLCELL_X1 FILLER_118_595 ();
 FILLCELL_X8 FILLER_118_600 ();
 FILLCELL_X1 FILLER_118_608 ();
 FILLCELL_X4 FILLER_118_632 ();
 FILLCELL_X1 FILLER_118_636 ();
 FILLCELL_X2 FILLER_118_648 ();
 FILLCELL_X2 FILLER_118_660 ();
 FILLCELL_X1 FILLER_118_676 ();
 FILLCELL_X1 FILLER_118_679 ();
 FILLCELL_X4 FILLER_118_705 ();
 FILLCELL_X2 FILLER_118_709 ();
 FILLCELL_X1 FILLER_118_711 ();
 FILLCELL_X8 FILLER_118_734 ();
 FILLCELL_X1 FILLER_118_742 ();
 FILLCELL_X16 FILLER_118_760 ();
 FILLCELL_X1 FILLER_118_776 ();
 FILLCELL_X2 FILLER_118_870 ();
 FILLCELL_X1 FILLER_118_872 ();
 FILLCELL_X1 FILLER_118_882 ();
 FILLCELL_X2 FILLER_118_895 ();
 FILLCELL_X8 FILLER_118_928 ();
 FILLCELL_X1 FILLER_118_936 ();
 FILLCELL_X2 FILLER_118_1009 ();
 FILLCELL_X2 FILLER_118_1018 ();
 FILLCELL_X32 FILLER_118_1036 ();
 FILLCELL_X4 FILLER_118_1068 ();
 FILLCELL_X16 FILLER_118_1080 ();
 FILLCELL_X4 FILLER_118_1096 ();
 FILLCELL_X2 FILLER_118_1100 ();
 FILLCELL_X1 FILLER_118_1102 ();
 FILLCELL_X4 FILLER_118_1111 ();
 FILLCELL_X2 FILLER_118_1115 ();
 FILLCELL_X4 FILLER_118_1121 ();
 FILLCELL_X16 FILLER_118_1129 ();
 FILLCELL_X2 FILLER_118_1145 ();
 FILLCELL_X1 FILLER_118_1147 ();
 FILLCELL_X1 FILLER_119_65 ();
 FILLCELL_X4 FILLER_119_68 ();
 FILLCELL_X2 FILLER_119_72 ();
 FILLCELL_X1 FILLER_119_78 ();
 FILLCELL_X4 FILLER_119_133 ();
 FILLCELL_X2 FILLER_119_137 ();
 FILLCELL_X1 FILLER_119_139 ();
 FILLCELL_X4 FILLER_119_194 ();
 FILLCELL_X2 FILLER_119_198 ();
 FILLCELL_X1 FILLER_119_228 ();
 FILLCELL_X1 FILLER_119_242 ();
 FILLCELL_X1 FILLER_119_267 ();
 FILLCELL_X1 FILLER_119_303 ();
 FILLCELL_X1 FILLER_119_440 ();
 FILLCELL_X4 FILLER_119_467 ();
 FILLCELL_X2 FILLER_119_475 ();
 FILLCELL_X1 FILLER_119_477 ();
 FILLCELL_X1 FILLER_119_484 ();
 FILLCELL_X2 FILLER_119_515 ();
 FILLCELL_X1 FILLER_119_532 ();
 FILLCELL_X1 FILLER_119_561 ();
 FILLCELL_X2 FILLER_119_573 ();
 FILLCELL_X2 FILLER_119_586 ();
 FILLCELL_X8 FILLER_119_591 ();
 FILLCELL_X1 FILLER_119_599 ();
 FILLCELL_X8 FILLER_119_618 ();
 FILLCELL_X2 FILLER_119_626 ();
 FILLCELL_X1 FILLER_119_651 ();
 FILLCELL_X1 FILLER_119_682 ();
 FILLCELL_X2 FILLER_119_726 ();
 FILLCELL_X1 FILLER_119_734 ();
 FILLCELL_X1 FILLER_119_745 ();
 FILLCELL_X1 FILLER_119_761 ();
 FILLCELL_X8 FILLER_119_780 ();
 FILLCELL_X4 FILLER_119_788 ();
 FILLCELL_X1 FILLER_119_812 ();
 FILLCELL_X1 FILLER_119_815 ();
 FILLCELL_X1 FILLER_119_868 ();
 FILLCELL_X2 FILLER_119_909 ();
 FILLCELL_X1 FILLER_119_911 ();
 FILLCELL_X2 FILLER_119_940 ();
 FILLCELL_X1 FILLER_119_976 ();
 FILLCELL_X1 FILLER_119_981 ();
 FILLCELL_X2 FILLER_119_1003 ();
 FILLCELL_X1 FILLER_119_1005 ();
 FILLCELL_X8 FILLER_119_1030 ();
 FILLCELL_X2 FILLER_119_1038 ();
 FILLCELL_X32 FILLER_119_1062 ();
 FILLCELL_X1 FILLER_119_1094 ();
 FILLCELL_X8 FILLER_119_1117 ();
 FILLCELL_X2 FILLER_119_1125 ();
 FILLCELL_X1 FILLER_119_1127 ();
 FILLCELL_X1 FILLER_120_1 ();
 FILLCELL_X1 FILLER_120_4 ();
 FILLCELL_X4 FILLER_120_37 ();
 FILLCELL_X2 FILLER_120_41 ();
 FILLCELL_X1 FILLER_120_51 ();
 FILLCELL_X2 FILLER_120_70 ();
 FILLCELL_X1 FILLER_120_72 ();
 FILLCELL_X8 FILLER_120_76 ();
 FILLCELL_X1 FILLER_120_87 ();
 FILLCELL_X8 FILLER_120_91 ();
 FILLCELL_X2 FILLER_120_99 ();
 FILLCELL_X1 FILLER_120_135 ();
 FILLCELL_X8 FILLER_120_138 ();
 FILLCELL_X1 FILLER_120_146 ();
 FILLCELL_X16 FILLER_120_151 ();
 FILLCELL_X1 FILLER_120_167 ();
 FILLCELL_X2 FILLER_120_193 ();
 FILLCELL_X1 FILLER_120_195 ();
 FILLCELL_X1 FILLER_120_209 ();
 FILLCELL_X1 FILLER_120_225 ();
 FILLCELL_X2 FILLER_120_247 ();
 FILLCELL_X1 FILLER_120_249 ();
 FILLCELL_X4 FILLER_120_271 ();
 FILLCELL_X2 FILLER_120_275 ();
 FILLCELL_X1 FILLER_120_277 ();
 FILLCELL_X1 FILLER_120_300 ();
 FILLCELL_X1 FILLER_120_309 ();
 FILLCELL_X1 FILLER_120_326 ();
 FILLCELL_X1 FILLER_120_374 ();
 FILLCELL_X1 FILLER_120_394 ();
 FILLCELL_X2 FILLER_120_411 ();
 FILLCELL_X1 FILLER_120_417 ();
 FILLCELL_X1 FILLER_120_429 ();
 FILLCELL_X1 FILLER_120_432 ();
 FILLCELL_X1 FILLER_120_463 ();
 FILLCELL_X2 FILLER_120_497 ();
 FILLCELL_X1 FILLER_120_499 ();
 FILLCELL_X2 FILLER_120_517 ();
 FILLCELL_X1 FILLER_120_519 ();
 FILLCELL_X1 FILLER_120_523 ();
 FILLCELL_X1 FILLER_120_529 ();
 FILLCELL_X2 FILLER_120_552 ();
 FILLCELL_X1 FILLER_120_559 ();
 FILLCELL_X1 FILLER_120_563 ();
 FILLCELL_X1 FILLER_120_575 ();
 FILLCELL_X2 FILLER_120_580 ();
 FILLCELL_X4 FILLER_120_600 ();
 FILLCELL_X2 FILLER_120_604 ();
 FILLCELL_X1 FILLER_120_606 ();
 FILLCELL_X4 FILLER_120_609 ();
 FILLCELL_X1 FILLER_120_613 ();
 FILLCELL_X1 FILLER_120_627 ();
 FILLCELL_X1 FILLER_120_630 ();
 FILLCELL_X1 FILLER_120_646 ();
 FILLCELL_X1 FILLER_120_700 ();
 FILLCELL_X1 FILLER_120_704 ();
 FILLCELL_X1 FILLER_120_712 ();
 FILLCELL_X1 FILLER_120_716 ();
 FILLCELL_X1 FILLER_120_722 ();
 FILLCELL_X1 FILLER_120_733 ();
 FILLCELL_X1 FILLER_120_767 ();
 FILLCELL_X2 FILLER_120_772 ();
 FILLCELL_X1 FILLER_120_774 ();
 FILLCELL_X1 FILLER_120_779 ();
 FILLCELL_X1 FILLER_120_782 ();
 FILLCELL_X2 FILLER_120_793 ();
 FILLCELL_X2 FILLER_120_800 ();
 FILLCELL_X1 FILLER_120_802 ();
 FILLCELL_X4 FILLER_120_838 ();
 FILLCELL_X1 FILLER_120_848 ();
 FILLCELL_X1 FILLER_120_852 ();
 FILLCELL_X4 FILLER_120_857 ();
 FILLCELL_X2 FILLER_120_861 ();
 FILLCELL_X1 FILLER_120_863 ();
 FILLCELL_X1 FILLER_120_873 ();
 FILLCELL_X1 FILLER_120_879 ();
 FILLCELL_X4 FILLER_120_900 ();
 FILLCELL_X2 FILLER_120_904 ();
 FILLCELL_X2 FILLER_120_913 ();
 FILLCELL_X1 FILLER_120_915 ();
 FILLCELL_X2 FILLER_120_945 ();
 FILLCELL_X1 FILLER_120_989 ();
 FILLCELL_X1 FILLER_120_999 ();
 FILLCELL_X1 FILLER_120_1007 ();
 FILLCELL_X32 FILLER_120_1044 ();
 FILLCELL_X32 FILLER_120_1076 ();
 FILLCELL_X16 FILLER_120_1108 ();
 FILLCELL_X4 FILLER_120_1124 ();
 FILLCELL_X1 FILLER_121_24 ();
 FILLCELL_X2 FILLER_121_97 ();
 FILLCELL_X1 FILLER_121_99 ();
 FILLCELL_X1 FILLER_121_139 ();
 FILLCELL_X1 FILLER_121_156 ();
 FILLCELL_X1 FILLER_121_177 ();
 FILLCELL_X2 FILLER_121_198 ();
 FILLCELL_X8 FILLER_121_214 ();
 FILLCELL_X1 FILLER_121_222 ();
 FILLCELL_X2 FILLER_121_258 ();
 FILLCELL_X1 FILLER_121_260 ();
 FILLCELL_X1 FILLER_121_287 ();
 FILLCELL_X1 FILLER_121_312 ();
 FILLCELL_X1 FILLER_121_323 ();
 FILLCELL_X2 FILLER_121_349 ();
 FILLCELL_X1 FILLER_121_387 ();
 FILLCELL_X2 FILLER_121_399 ();
 FILLCELL_X2 FILLER_121_465 ();
 FILLCELL_X1 FILLER_121_470 ();
 FILLCELL_X1 FILLER_121_502 ();
 FILLCELL_X1 FILLER_121_512 ();
 FILLCELL_X1 FILLER_121_538 ();
 FILLCELL_X4 FILLER_121_541 ();
 FILLCELL_X2 FILLER_121_552 ();
 FILLCELL_X1 FILLER_121_554 ();
 FILLCELL_X2 FILLER_121_565 ();
 FILLCELL_X1 FILLER_121_570 ();
 FILLCELL_X2 FILLER_121_616 ();
 FILLCELL_X1 FILLER_121_618 ();
 FILLCELL_X1 FILLER_121_632 ();
 FILLCELL_X2 FILLER_121_717 ();
 FILLCELL_X2 FILLER_121_726 ();
 FILLCELL_X1 FILLER_121_738 ();
 FILLCELL_X1 FILLER_121_743 ();
 FILLCELL_X1 FILLER_121_766 ();
 FILLCELL_X2 FILLER_121_777 ();
 FILLCELL_X2 FILLER_121_817 ();
 FILLCELL_X1 FILLER_121_838 ();
 FILLCELL_X1 FILLER_121_845 ();
 FILLCELL_X8 FILLER_121_862 ();
 FILLCELL_X16 FILLER_121_876 ();
 FILLCELL_X8 FILLER_121_892 ();
 FILLCELL_X2 FILLER_121_900 ();
 FILLCELL_X16 FILLER_121_950 ();
 FILLCELL_X8 FILLER_121_966 ();
 FILLCELL_X1 FILLER_121_974 ();
 FILLCELL_X8 FILLER_121_995 ();
 FILLCELL_X1 FILLER_121_1003 ();
 FILLCELL_X1 FILLER_121_1011 ();
 FILLCELL_X2 FILLER_121_1037 ();
 FILLCELL_X1 FILLER_121_1039 ();
 FILLCELL_X32 FILLER_121_1070 ();
 FILLCELL_X16 FILLER_121_1102 ();
 FILLCELL_X4 FILLER_121_1118 ();
 FILLCELL_X2 FILLER_121_1122 ();
 FILLCELL_X16 FILLER_121_1132 ();
 FILLCELL_X4 FILLER_122_25 ();
 FILLCELL_X1 FILLER_122_29 ();
 FILLCELL_X1 FILLER_122_42 ();
 FILLCELL_X4 FILLER_122_45 ();
 FILLCELL_X1 FILLER_122_53 ();
 FILLCELL_X1 FILLER_122_84 ();
 FILLCELL_X2 FILLER_122_87 ();
 FILLCELL_X8 FILLER_122_92 ();
 FILLCELL_X4 FILLER_122_100 ();
 FILLCELL_X1 FILLER_122_123 ();
 FILLCELL_X1 FILLER_122_160 ();
 FILLCELL_X2 FILLER_122_163 ();
 FILLCELL_X8 FILLER_122_169 ();
 FILLCELL_X2 FILLER_122_177 ();
 FILLCELL_X2 FILLER_122_278 ();
 FILLCELL_X4 FILLER_122_374 ();
 FILLCELL_X2 FILLER_122_378 ();
 FILLCELL_X1 FILLER_122_452 ();
 FILLCELL_X2 FILLER_122_473 ();
 FILLCELL_X2 FILLER_122_518 ();
 FILLCELL_X1 FILLER_122_528 ();
 FILLCELL_X1 FILLER_122_536 ();
 FILLCELL_X4 FILLER_122_575 ();
 FILLCELL_X4 FILLER_122_601 ();
 FILLCELL_X1 FILLER_122_605 ();
 FILLCELL_X2 FILLER_122_608 ();
 FILLCELL_X1 FILLER_122_610 ();
 FILLCELL_X2 FILLER_122_638 ();
 FILLCELL_X1 FILLER_122_640 ();
 FILLCELL_X2 FILLER_122_652 ();
 FILLCELL_X1 FILLER_122_669 ();
 FILLCELL_X2 FILLER_122_727 ();
 FILLCELL_X1 FILLER_122_783 ();
 FILLCELL_X2 FILLER_122_790 ();
 FILLCELL_X1 FILLER_122_792 ();
 FILLCELL_X16 FILLER_122_795 ();
 FILLCELL_X8 FILLER_122_811 ();
 FILLCELL_X2 FILLER_122_819 ();
 FILLCELL_X1 FILLER_122_821 ();
 FILLCELL_X2 FILLER_122_829 ();
 FILLCELL_X1 FILLER_122_831 ();
 FILLCELL_X1 FILLER_122_846 ();
 FILLCELL_X1 FILLER_122_849 ();
 FILLCELL_X1 FILLER_122_852 ();
 FILLCELL_X2 FILLER_122_867 ();
 FILLCELL_X1 FILLER_122_869 ();
 FILLCELL_X4 FILLER_122_883 ();
 FILLCELL_X2 FILLER_122_887 ();
 FILLCELL_X4 FILLER_122_909 ();
 FILLCELL_X2 FILLER_122_913 ();
 FILLCELL_X1 FILLER_122_915 ();
 FILLCELL_X1 FILLER_122_933 ();
 FILLCELL_X2 FILLER_122_948 ();
 FILLCELL_X1 FILLER_122_950 ();
 FILLCELL_X1 FILLER_122_967 ();
 FILLCELL_X16 FILLER_122_992 ();
 FILLCELL_X8 FILLER_122_1008 ();
 FILLCELL_X2 FILLER_122_1016 ();
 FILLCELL_X1 FILLER_122_1018 ();
 FILLCELL_X8 FILLER_122_1021 ();
 FILLCELL_X1 FILLER_122_1029 ();
 FILLCELL_X1 FILLER_122_1041 ();
 FILLCELL_X2 FILLER_122_1052 ();
 FILLCELL_X1 FILLER_122_1054 ();
 FILLCELL_X32 FILLER_122_1067 ();
 FILLCELL_X16 FILLER_122_1099 ();
 FILLCELL_X1 FILLER_122_1115 ();
 FILLCELL_X8 FILLER_122_1136 ();
 FILLCELL_X4 FILLER_122_1144 ();
 FILLCELL_X1 FILLER_123_15 ();
 FILLCELL_X2 FILLER_123_32 ();
 FILLCELL_X2 FILLER_123_37 ();
 FILLCELL_X2 FILLER_123_48 ();
 FILLCELL_X1 FILLER_123_50 ();
 FILLCELL_X2 FILLER_123_63 ();
 FILLCELL_X1 FILLER_123_68 ();
 FILLCELL_X2 FILLER_123_101 ();
 FILLCELL_X2 FILLER_123_108 ();
 FILLCELL_X1 FILLER_123_110 ();
 FILLCELL_X2 FILLER_123_181 ();
 FILLCELL_X1 FILLER_123_183 ();
 FILLCELL_X4 FILLER_123_208 ();
 FILLCELL_X2 FILLER_123_244 ();
 FILLCELL_X2 FILLER_123_254 ();
 FILLCELL_X1 FILLER_123_306 ();
 FILLCELL_X2 FILLER_123_367 ();
 FILLCELL_X4 FILLER_123_394 ();
 FILLCELL_X1 FILLER_123_428 ();
 FILLCELL_X1 FILLER_123_480 ();
 FILLCELL_X1 FILLER_123_484 ();
 FILLCELL_X2 FILLER_123_495 ();
 FILLCELL_X2 FILLER_123_507 ();
 FILLCELL_X2 FILLER_123_519 ();
 FILLCELL_X1 FILLER_123_521 ();
 FILLCELL_X1 FILLER_123_536 ();
 FILLCELL_X1 FILLER_123_541 ();
 FILLCELL_X1 FILLER_123_544 ();
 FILLCELL_X4 FILLER_123_557 ();
 FILLCELL_X4 FILLER_123_563 ();
 FILLCELL_X2 FILLER_123_567 ();
 FILLCELL_X1 FILLER_123_569 ();
 FILLCELL_X4 FILLER_123_588 ();
 FILLCELL_X1 FILLER_123_592 ();
 FILLCELL_X2 FILLER_123_595 ();
 FILLCELL_X1 FILLER_123_597 ();
 FILLCELL_X4 FILLER_123_638 ();
 FILLCELL_X2 FILLER_123_652 ();
 FILLCELL_X2 FILLER_123_680 ();
 FILLCELL_X2 FILLER_123_726 ();
 FILLCELL_X4 FILLER_123_759 ();
 FILLCELL_X2 FILLER_123_763 ();
 FILLCELL_X8 FILLER_123_806 ();
 FILLCELL_X2 FILLER_123_814 ();
 FILLCELL_X1 FILLER_123_840 ();
 FILLCELL_X8 FILLER_123_857 ();
 FILLCELL_X2 FILLER_123_916 ();
 FILLCELL_X1 FILLER_123_918 ();
 FILLCELL_X8 FILLER_123_934 ();
 FILLCELL_X1 FILLER_123_942 ();
 FILLCELL_X2 FILLER_123_950 ();
 FILLCELL_X1 FILLER_123_952 ();
 FILLCELL_X8 FILLER_123_1002 ();
 FILLCELL_X4 FILLER_123_1010 ();
 FILLCELL_X2 FILLER_123_1019 ();
 FILLCELL_X2 FILLER_123_1028 ();
 FILLCELL_X2 FILLER_123_1040 ();
 FILLCELL_X1 FILLER_123_1042 ();
 FILLCELL_X1 FILLER_123_1045 ();
 FILLCELL_X2 FILLER_123_1050 ();
 FILLCELL_X1 FILLER_123_1052 ();
 FILLCELL_X8 FILLER_123_1067 ();
 FILLCELL_X4 FILLER_123_1075 ();
 FILLCELL_X32 FILLER_123_1091 ();
 FILLCELL_X2 FILLER_123_1123 ();
 FILLCELL_X2 FILLER_123_1145 ();
 FILLCELL_X1 FILLER_123_1147 ();
 FILLCELL_X1 FILLER_124_1 ();
 FILLCELL_X2 FILLER_124_46 ();
 FILLCELL_X2 FILLER_124_60 ();
 FILLCELL_X8 FILLER_124_76 ();
 FILLCELL_X4 FILLER_124_84 ();
 FILLCELL_X2 FILLER_124_88 ();
 FILLCELL_X1 FILLER_124_90 ();
 FILLCELL_X8 FILLER_124_127 ();
 FILLCELL_X2 FILLER_124_135 ();
 FILLCELL_X1 FILLER_124_137 ();
 FILLCELL_X16 FILLER_124_140 ();
 FILLCELL_X2 FILLER_124_156 ();
 FILLCELL_X2 FILLER_124_161 ();
 FILLCELL_X8 FILLER_124_168 ();
 FILLCELL_X2 FILLER_124_176 ();
 FILLCELL_X2 FILLER_124_213 ();
 FILLCELL_X1 FILLER_124_215 ();
 FILLCELL_X8 FILLER_124_226 ();
 FILLCELL_X2 FILLER_124_234 ();
 FILLCELL_X8 FILLER_124_288 ();
 FILLCELL_X2 FILLER_124_338 ();
 FILLCELL_X8 FILLER_124_402 ();
 FILLCELL_X2 FILLER_124_410 ();
 FILLCELL_X1 FILLER_124_412 ();
 FILLCELL_X1 FILLER_124_433 ();
 FILLCELL_X2 FILLER_124_464 ();
 FILLCELL_X1 FILLER_124_479 ();
 FILLCELL_X1 FILLER_124_528 ();
 FILLCELL_X2 FILLER_124_549 ();
 FILLCELL_X2 FILLER_124_569 ();
 FILLCELL_X8 FILLER_124_587 ();
 FILLCELL_X2 FILLER_124_597 ();
 FILLCELL_X4 FILLER_124_624 ();
 FILLCELL_X2 FILLER_124_628 ();
 FILLCELL_X1 FILLER_124_630 ();
 FILLCELL_X4 FILLER_124_714 ();
 FILLCELL_X1 FILLER_124_728 ();
 FILLCELL_X2 FILLER_124_749 ();
 FILLCELL_X2 FILLER_124_771 ();
 FILLCELL_X2 FILLER_124_793 ();
 FILLCELL_X16 FILLER_124_805 ();
 FILLCELL_X2 FILLER_124_821 ();
 FILLCELL_X2 FILLER_124_831 ();
 FILLCELL_X1 FILLER_124_833 ();
 FILLCELL_X1 FILLER_124_864 ();
 FILLCELL_X2 FILLER_124_901 ();
 FILLCELL_X2 FILLER_124_913 ();
 FILLCELL_X1 FILLER_124_929 ();
 FILLCELL_X4 FILLER_124_935 ();
 FILLCELL_X2 FILLER_124_939 ();
 FILLCELL_X1 FILLER_124_941 ();
 FILLCELL_X8 FILLER_124_946 ();
 FILLCELL_X4 FILLER_124_954 ();
 FILLCELL_X1 FILLER_124_958 ();
 FILLCELL_X2 FILLER_124_1018 ();
 FILLCELL_X1 FILLER_124_1063 ();
 FILLCELL_X2 FILLER_124_1071 ();
 FILLCELL_X1 FILLER_124_1073 ();
 FILLCELL_X8 FILLER_124_1092 ();
 FILLCELL_X2 FILLER_124_1100 ();
 FILLCELL_X16 FILLER_124_1122 ();
 FILLCELL_X4 FILLER_124_1138 ();
 FILLCELL_X2 FILLER_124_1142 ();
 FILLCELL_X1 FILLER_124_1144 ();
 FILLCELL_X2 FILLER_125_4 ();
 FILLCELL_X2 FILLER_125_12 ();
 FILLCELL_X1 FILLER_125_26 ();
 FILLCELL_X1 FILLER_125_45 ();
 FILLCELL_X1 FILLER_125_62 ();
 FILLCELL_X1 FILLER_125_81 ();
 FILLCELL_X4 FILLER_125_84 ();
 FILLCELL_X2 FILLER_125_88 ();
 FILLCELL_X1 FILLER_125_92 ();
 FILLCELL_X8 FILLER_125_105 ();
 FILLCELL_X2 FILLER_125_113 ();
 FILLCELL_X4 FILLER_125_119 ();
 FILLCELL_X2 FILLER_125_123 ();
 FILLCELL_X1 FILLER_125_125 ();
 FILLCELL_X2 FILLER_125_136 ();
 FILLCELL_X1 FILLER_125_138 ();
 FILLCELL_X2 FILLER_125_149 ();
 FILLCELL_X1 FILLER_125_151 ();
 FILLCELL_X2 FILLER_125_170 ();
 FILLCELL_X2 FILLER_125_188 ();
 FILLCELL_X8 FILLER_125_194 ();
 FILLCELL_X2 FILLER_125_202 ();
 FILLCELL_X4 FILLER_125_208 ();
 FILLCELL_X2 FILLER_125_212 ();
 FILLCELL_X4 FILLER_125_236 ();
 FILLCELL_X2 FILLER_125_240 ();
 FILLCELL_X1 FILLER_125_262 ();
 FILLCELL_X4 FILLER_125_268 ();
 FILLCELL_X2 FILLER_125_272 ();
 FILLCELL_X16 FILLER_125_276 ();
 FILLCELL_X4 FILLER_125_292 ();
 FILLCELL_X1 FILLER_125_300 ();
 FILLCELL_X1 FILLER_125_305 ();
 FILLCELL_X2 FILLER_125_310 ();
 FILLCELL_X2 FILLER_125_318 ();
 FILLCELL_X2 FILLER_125_336 ();
 FILLCELL_X4 FILLER_125_340 ();
 FILLCELL_X1 FILLER_125_344 ();
 FILLCELL_X16 FILLER_125_347 ();
 FILLCELL_X8 FILLER_125_363 ();
 FILLCELL_X4 FILLER_125_371 ();
 FILLCELL_X2 FILLER_125_388 ();
 FILLCELL_X2 FILLER_125_392 ();
 FILLCELL_X2 FILLER_125_434 ();
 FILLCELL_X4 FILLER_125_445 ();
 FILLCELL_X4 FILLER_125_534 ();
 FILLCELL_X1 FILLER_125_538 ();
 FILLCELL_X8 FILLER_125_547 ();
 FILLCELL_X2 FILLER_125_571 ();
 FILLCELL_X2 FILLER_125_577 ();
 FILLCELL_X1 FILLER_125_579 ();
 FILLCELL_X8 FILLER_125_596 ();
 FILLCELL_X2 FILLER_125_604 ();
 FILLCELL_X1 FILLER_125_606 ();
 FILLCELL_X8 FILLER_125_609 ();
 FILLCELL_X1 FILLER_125_619 ();
 FILLCELL_X8 FILLER_125_650 ();
 FILLCELL_X4 FILLER_125_684 ();
 FILLCELL_X8 FILLER_125_693 ();
 FILLCELL_X2 FILLER_125_701 ();
 FILLCELL_X1 FILLER_125_723 ();
 FILLCELL_X8 FILLER_125_744 ();
 FILLCELL_X1 FILLER_125_752 ();
 FILLCELL_X4 FILLER_125_773 ();
 FILLCELL_X2 FILLER_125_777 ();
 FILLCELL_X1 FILLER_125_779 ();
 FILLCELL_X2 FILLER_125_850 ();
 FILLCELL_X1 FILLER_125_858 ();
 FILLCELL_X1 FILLER_125_865 ();
 FILLCELL_X4 FILLER_125_878 ();
 FILLCELL_X2 FILLER_125_882 ();
 FILLCELL_X1 FILLER_125_904 ();
 FILLCELL_X2 FILLER_125_932 ();
 FILLCELL_X2 FILLER_125_946 ();
 FILLCELL_X1 FILLER_125_948 ();
 FILLCELL_X8 FILLER_125_954 ();
 FILLCELL_X1 FILLER_125_962 ();
 FILLCELL_X4 FILLER_125_977 ();
 FILLCELL_X1 FILLER_125_981 ();
 FILLCELL_X4 FILLER_125_989 ();
 FILLCELL_X1 FILLER_125_993 ();
 FILLCELL_X1 FILLER_125_1001 ();
 FILLCELL_X2 FILLER_125_1016 ();
 FILLCELL_X8 FILLER_125_1025 ();
 FILLCELL_X2 FILLER_125_1080 ();
 FILLCELL_X8 FILLER_125_1110 ();
 FILLCELL_X4 FILLER_125_1118 ();
 FILLCELL_X1 FILLER_125_1122 ();
 FILLCELL_X2 FILLER_125_1143 ();
 FILLCELL_X1 FILLER_126_17 ();
 FILLCELL_X2 FILLER_126_34 ();
 FILLCELL_X1 FILLER_126_36 ();
 FILLCELL_X2 FILLER_126_41 ();
 FILLCELL_X2 FILLER_126_51 ();
 FILLCELL_X4 FILLER_126_57 ();
 FILLCELL_X2 FILLER_126_61 ();
 FILLCELL_X1 FILLER_126_63 ();
 FILLCELL_X1 FILLER_126_66 ();
 FILLCELL_X2 FILLER_126_69 ();
 FILLCELL_X1 FILLER_126_115 ();
 FILLCELL_X1 FILLER_126_120 ();
 FILLCELL_X1 FILLER_126_137 ();
 FILLCELL_X1 FILLER_126_154 ();
 FILLCELL_X1 FILLER_126_166 ();
 FILLCELL_X2 FILLER_126_204 ();
 FILLCELL_X1 FILLER_126_206 ();
 FILLCELL_X2 FILLER_126_223 ();
 FILLCELL_X8 FILLER_126_255 ();
 FILLCELL_X2 FILLER_126_263 ();
 FILLCELL_X8 FILLER_126_275 ();
 FILLCELL_X4 FILLER_126_283 ();
 FILLCELL_X2 FILLER_126_287 ();
 FILLCELL_X1 FILLER_126_289 ();
 FILLCELL_X2 FILLER_126_306 ();
 FILLCELL_X1 FILLER_126_310 ();
 FILLCELL_X8 FILLER_126_313 ();
 FILLCELL_X4 FILLER_126_321 ();
 FILLCELL_X2 FILLER_126_325 ();
 FILLCELL_X1 FILLER_126_327 ();
 FILLCELL_X4 FILLER_126_330 ();
 FILLCELL_X2 FILLER_126_334 ();
 FILLCELL_X1 FILLER_126_336 ();
 FILLCELL_X1 FILLER_126_364 ();
 FILLCELL_X8 FILLER_126_385 ();
 FILLCELL_X4 FILLER_126_393 ();
 FILLCELL_X1 FILLER_126_413 ();
 FILLCELL_X8 FILLER_126_418 ();
 FILLCELL_X4 FILLER_126_426 ();
 FILLCELL_X4 FILLER_126_472 ();
 FILLCELL_X8 FILLER_126_501 ();
 FILLCELL_X4 FILLER_126_509 ();
 FILLCELL_X1 FILLER_126_513 ();
 FILLCELL_X4 FILLER_126_516 ();
 FILLCELL_X1 FILLER_126_520 ();
 FILLCELL_X2 FILLER_126_551 ();
 FILLCELL_X2 FILLER_126_563 ();
 FILLCELL_X1 FILLER_126_565 ();
 FILLCELL_X4 FILLER_126_569 ();
 FILLCELL_X1 FILLER_126_573 ();
 FILLCELL_X1 FILLER_126_580 ();
 FILLCELL_X4 FILLER_126_585 ();
 FILLCELL_X4 FILLER_126_592 ();
 FILLCELL_X1 FILLER_126_596 ();
 FILLCELL_X2 FILLER_126_599 ();
 FILLCELL_X8 FILLER_126_623 ();
 FILLCELL_X1 FILLER_126_632 ();
 FILLCELL_X16 FILLER_126_675 ();
 FILLCELL_X8 FILLER_126_691 ();
 FILLCELL_X1 FILLER_126_699 ();
 FILLCELL_X2 FILLER_126_722 ();
 FILLCELL_X1 FILLER_126_724 ();
 FILLCELL_X4 FILLER_126_749 ();
 FILLCELL_X2 FILLER_126_753 ();
 FILLCELL_X4 FILLER_126_760 ();
 FILLCELL_X2 FILLER_126_764 ();
 FILLCELL_X1 FILLER_126_766 ();
 FILLCELL_X4 FILLER_126_797 ();
 FILLCELL_X2 FILLER_126_801 ();
 FILLCELL_X1 FILLER_126_803 ();
 FILLCELL_X8 FILLER_126_824 ();
 FILLCELL_X4 FILLER_126_832 ();
 FILLCELL_X2 FILLER_126_836 ();
 FILLCELL_X1 FILLER_126_838 ();
 FILLCELL_X1 FILLER_126_859 ();
 FILLCELL_X1 FILLER_126_925 ();
 FILLCELL_X4 FILLER_126_930 ();
 FILLCELL_X2 FILLER_126_934 ();
 FILLCELL_X1 FILLER_126_936 ();
 FILLCELL_X4 FILLER_126_945 ();
 FILLCELL_X2 FILLER_126_949 ();
 FILLCELL_X1 FILLER_126_951 ();
 FILLCELL_X1 FILLER_126_1009 ();
 FILLCELL_X1 FILLER_126_1016 ();
 FILLCELL_X1 FILLER_126_1019 ();
 FILLCELL_X1 FILLER_126_1036 ();
 FILLCELL_X4 FILLER_126_1053 ();
 FILLCELL_X1 FILLER_126_1057 ();
 FILLCELL_X1 FILLER_126_1093 ();
 FILLCELL_X1 FILLER_126_1098 ();
 FILLCELL_X1 FILLER_126_1108 ();
 FILLCELL_X1 FILLER_126_1116 ();
 FILLCELL_X1 FILLER_126_1144 ();
 FILLCELL_X1 FILLER_127_1 ();
 FILLCELL_X1 FILLER_127_9 ();
 FILLCELL_X8 FILLER_127_26 ();
 FILLCELL_X1 FILLER_127_34 ();
 FILLCELL_X1 FILLER_127_57 ();
 FILLCELL_X4 FILLER_127_74 ();
 FILLCELL_X2 FILLER_127_78 ();
 FILLCELL_X1 FILLER_127_80 ();
 FILLCELL_X2 FILLER_127_83 ();
 FILLCELL_X4 FILLER_127_87 ();
 FILLCELL_X8 FILLER_127_119 ();
 FILLCELL_X8 FILLER_127_131 ();
 FILLCELL_X2 FILLER_127_167 ();
 FILLCELL_X2 FILLER_127_185 ();
 FILLCELL_X1 FILLER_127_203 ();
 FILLCELL_X2 FILLER_127_218 ();
 FILLCELL_X8 FILLER_127_245 ();
 FILLCELL_X4 FILLER_127_280 ();
 FILLCELL_X2 FILLER_127_284 ();
 FILLCELL_X1 FILLER_127_286 ();
 FILLCELL_X1 FILLER_127_291 ();
 FILLCELL_X1 FILLER_127_296 ();
 FILLCELL_X1 FILLER_127_317 ();
 FILLCELL_X8 FILLER_127_365 ();
 FILLCELL_X8 FILLER_127_405 ();
 FILLCELL_X2 FILLER_127_413 ();
 FILLCELL_X1 FILLER_127_431 ();
 FILLCELL_X1 FILLER_127_450 ();
 FILLCELL_X1 FILLER_127_453 ();
 FILLCELL_X8 FILLER_127_456 ();
 FILLCELL_X4 FILLER_127_464 ();
 FILLCELL_X2 FILLER_127_492 ();
 FILLCELL_X8 FILLER_127_514 ();
 FILLCELL_X4 FILLER_127_546 ();
 FILLCELL_X1 FILLER_127_602 ();
 FILLCELL_X8 FILLER_127_626 ();
 FILLCELL_X8 FILLER_127_658 ();
 FILLCELL_X4 FILLER_127_666 ();
 FILLCELL_X8 FILLER_127_672 ();
 FILLCELL_X1 FILLER_127_682 ();
 FILLCELL_X2 FILLER_127_701 ();
 FILLCELL_X1 FILLER_127_703 ();
 FILLCELL_X8 FILLER_127_706 ();
 FILLCELL_X1 FILLER_127_714 ();
 FILLCELL_X2 FILLER_127_735 ();
 FILLCELL_X1 FILLER_127_737 ();
 FILLCELL_X2 FILLER_127_758 ();
 FILLCELL_X4 FILLER_127_770 ();
 FILLCELL_X2 FILLER_127_774 ();
 FILLCELL_X1 FILLER_127_776 ();
 FILLCELL_X4 FILLER_127_781 ();
 FILLCELL_X4 FILLER_127_805 ();
 FILLCELL_X2 FILLER_127_809 ();
 FILLCELL_X1 FILLER_127_811 ();
 FILLCELL_X1 FILLER_127_834 ();
 FILLCELL_X4 FILLER_127_856 ();
 FILLCELL_X2 FILLER_127_860 ();
 FILLCELL_X1 FILLER_127_862 ();
 FILLCELL_X2 FILLER_127_883 ();
 FILLCELL_X1 FILLER_127_885 ();
 FILLCELL_X2 FILLER_127_934 ();
 FILLCELL_X8 FILLER_127_956 ();
 FILLCELL_X2 FILLER_127_964 ();
 FILLCELL_X1 FILLER_127_1009 ();
 FILLCELL_X1 FILLER_127_1051 ();
 FILLCELL_X2 FILLER_127_1146 ();
 FILLCELL_X1 FILLER_128_1 ();
 FILLCELL_X2 FILLER_128_45 ();
 FILLCELL_X1 FILLER_128_47 ();
 FILLCELL_X2 FILLER_128_52 ();
 FILLCELL_X1 FILLER_128_54 ();
 FILLCELL_X2 FILLER_128_57 ();
 FILLCELL_X1 FILLER_128_59 ();
 FILLCELL_X4 FILLER_128_62 ();
 FILLCELL_X2 FILLER_128_66 ();
 FILLCELL_X2 FILLER_128_131 ();
 FILLCELL_X1 FILLER_128_133 ();
 FILLCELL_X2 FILLER_128_140 ();
 FILLCELL_X1 FILLER_128_142 ();
 FILLCELL_X1 FILLER_128_155 ();
 FILLCELL_X1 FILLER_128_164 ();
 FILLCELL_X1 FILLER_128_181 ();
 FILLCELL_X2 FILLER_128_191 ();
 FILLCELL_X1 FILLER_128_193 ();
 FILLCELL_X2 FILLER_128_202 ();
 FILLCELL_X2 FILLER_128_215 ();
 FILLCELL_X8 FILLER_128_257 ();
 FILLCELL_X4 FILLER_128_265 ();
 FILLCELL_X2 FILLER_128_269 ();
 FILLCELL_X1 FILLER_128_271 ();
 FILLCELL_X2 FILLER_128_290 ();
 FILLCELL_X1 FILLER_128_292 ();
 FILLCELL_X2 FILLER_128_304 ();
 FILLCELL_X1 FILLER_128_306 ();
 FILLCELL_X4 FILLER_128_309 ();
 FILLCELL_X1 FILLER_128_329 ();
 FILLCELL_X1 FILLER_128_346 ();
 FILLCELL_X8 FILLER_128_349 ();
 FILLCELL_X4 FILLER_128_389 ();
 FILLCELL_X2 FILLER_128_395 ();
 FILLCELL_X1 FILLER_128_399 ();
 FILLCELL_X1 FILLER_128_403 ();
 FILLCELL_X2 FILLER_128_422 ();
 FILLCELL_X1 FILLER_128_424 ();
 FILLCELL_X4 FILLER_128_441 ();
 FILLCELL_X1 FILLER_128_445 ();
 FILLCELL_X4 FILLER_128_448 ();
 FILLCELL_X1 FILLER_128_452 ();
 FILLCELL_X2 FILLER_128_469 ();
 FILLCELL_X1 FILLER_128_471 ();
 FILLCELL_X1 FILLER_128_474 ();
 FILLCELL_X1 FILLER_128_477 ();
 FILLCELL_X4 FILLER_128_496 ();
 FILLCELL_X2 FILLER_128_500 ();
 FILLCELL_X1 FILLER_128_502 ();
 FILLCELL_X1 FILLER_128_522 ();
 FILLCELL_X4 FILLER_128_530 ();
 FILLCELL_X2 FILLER_128_534 ();
 FILLCELL_X2 FILLER_128_552 ();
 FILLCELL_X1 FILLER_128_558 ();
 FILLCELL_X1 FILLER_128_579 ();
 FILLCELL_X2 FILLER_128_584 ();
 FILLCELL_X1 FILLER_128_586 ();
 FILLCELL_X1 FILLER_128_605 ();
 FILLCELL_X1 FILLER_128_635 ();
 FILLCELL_X2 FILLER_128_716 ();
 FILLCELL_X8 FILLER_128_720 ();
 FILLCELL_X2 FILLER_128_728 ();
 FILLCELL_X1 FILLER_128_784 ();
 FILLCELL_X4 FILLER_128_789 ();
 FILLCELL_X2 FILLER_128_793 ();
 FILLCELL_X4 FILLER_128_815 ();
 FILLCELL_X2 FILLER_128_819 ();
 FILLCELL_X1 FILLER_128_821 ();
 FILLCELL_X4 FILLER_128_853 ();
 FILLCELL_X1 FILLER_128_857 ();
 FILLCELL_X1 FILLER_128_878 ();
 FILLCELL_X1 FILLER_128_899 ();
 FILLCELL_X1 FILLER_128_903 ();
 FILLCELL_X1 FILLER_128_914 ();
 FILLCELL_X1 FILLER_128_920 ();
 FILLCELL_X1 FILLER_128_933 ();
 FILLCELL_X2 FILLER_128_971 ();
 FILLCELL_X1 FILLER_128_973 ();
 FILLCELL_X1 FILLER_128_981 ();
 FILLCELL_X1 FILLER_128_986 ();
 FILLCELL_X2 FILLER_128_991 ();
 FILLCELL_X4 FILLER_128_1020 ();
 FILLCELL_X1 FILLER_128_1089 ();
 FILLCELL_X1 FILLER_128_1099 ();
 FILLCELL_X1 FILLER_128_1123 ();
 FILLCELL_X1 FILLER_128_1147 ();
 FILLCELL_X1 FILLER_129_4 ();
 FILLCELL_X2 FILLER_129_13 ();
 FILLCELL_X2 FILLER_129_84 ();
 FILLCELL_X4 FILLER_129_108 ();
 FILLCELL_X2 FILLER_129_112 ();
 FILLCELL_X1 FILLER_129_114 ();
 FILLCELL_X4 FILLER_129_117 ();
 FILLCELL_X2 FILLER_129_121 ();
 FILLCELL_X1 FILLER_129_123 ();
 FILLCELL_X4 FILLER_129_144 ();
 FILLCELL_X1 FILLER_129_168 ();
 FILLCELL_X8 FILLER_129_219 ();
 FILLCELL_X4 FILLER_129_239 ();
 FILLCELL_X1 FILLER_129_243 ();
 FILLCELL_X4 FILLER_129_258 ();
 FILLCELL_X2 FILLER_129_288 ();
 FILLCELL_X1 FILLER_129_290 ();
 FILLCELL_X2 FILLER_129_343 ();
 FILLCELL_X1 FILLER_129_462 ();
 FILLCELL_X1 FILLER_129_466 ();
 FILLCELL_X1 FILLER_129_483 ();
 FILLCELL_X2 FILLER_129_486 ();
 FILLCELL_X16 FILLER_129_492 ();
 FILLCELL_X4 FILLER_129_508 ();
 FILLCELL_X1 FILLER_129_514 ();
 FILLCELL_X1 FILLER_129_518 ();
 FILLCELL_X2 FILLER_129_539 ();
 FILLCELL_X2 FILLER_129_558 ();
 FILLCELL_X1 FILLER_129_560 ();
 FILLCELL_X4 FILLER_129_599 ();
 FILLCELL_X2 FILLER_129_603 ();
 FILLCELL_X2 FILLER_129_607 ();
 FILLCELL_X4 FILLER_129_611 ();
 FILLCELL_X2 FILLER_129_643 ();
 FILLCELL_X1 FILLER_129_645 ();
 FILLCELL_X2 FILLER_129_662 ();
 FILLCELL_X1 FILLER_129_666 ();
 FILLCELL_X2 FILLER_129_671 ();
 FILLCELL_X1 FILLER_129_689 ();
 FILLCELL_X1 FILLER_129_692 ();
 FILLCELL_X1 FILLER_129_695 ();
 FILLCELL_X1 FILLER_129_699 ();
 FILLCELL_X4 FILLER_129_735 ();
 FILLCELL_X2 FILLER_129_741 ();
 FILLCELL_X4 FILLER_129_745 ();
 FILLCELL_X2 FILLER_129_749 ();
 FILLCELL_X1 FILLER_129_759 ();
 FILLCELL_X1 FILLER_129_764 ();
 FILLCELL_X2 FILLER_129_769 ();
 FILLCELL_X1 FILLER_129_779 ();
 FILLCELL_X4 FILLER_129_784 ();
 FILLCELL_X4 FILLER_129_808 ();
 FILLCELL_X2 FILLER_129_837 ();
 FILLCELL_X2 FILLER_129_848 ();
 FILLCELL_X1 FILLER_129_850 ();
 FILLCELL_X2 FILLER_129_878 ();
 FILLCELL_X1 FILLER_129_903 ();
 FILLCELL_X1 FILLER_129_910 ();
 FILLCELL_X1 FILLER_129_922 ();
 FILLCELL_X1 FILLER_129_926 ();
 FILLCELL_X4 FILLER_129_934 ();
 FILLCELL_X2 FILLER_129_938 ();
 FILLCELL_X1 FILLER_129_940 ();
 FILLCELL_X2 FILLER_129_951 ();
 FILLCELL_X1 FILLER_129_953 ();
 FILLCELL_X4 FILLER_129_957 ();
 FILLCELL_X1 FILLER_129_961 ();
 FILLCELL_X2 FILLER_129_976 ();
 FILLCELL_X1 FILLER_129_985 ();
 FILLCELL_X2 FILLER_129_993 ();
 FILLCELL_X2 FILLER_129_999 ();
 FILLCELL_X2 FILLER_129_1037 ();
 FILLCELL_X2 FILLER_129_1043 ();
 FILLCELL_X1 FILLER_129_1064 ();
 FILLCELL_X1 FILLER_129_1088 ();
 FILLCELL_X4 FILLER_130_1 ();
 FILLCELL_X2 FILLER_130_5 ();
 FILLCELL_X1 FILLER_130_7 ();
 FILLCELL_X4 FILLER_130_24 ();
 FILLCELL_X2 FILLER_130_28 ();
 FILLCELL_X1 FILLER_130_30 ();
 FILLCELL_X16 FILLER_130_87 ();
 FILLCELL_X4 FILLER_130_103 ();
 FILLCELL_X2 FILLER_130_107 ();
 FILLCELL_X2 FILLER_130_111 ();
 FILLCELL_X2 FILLER_130_135 ();
 FILLCELL_X1 FILLER_130_137 ();
 FILLCELL_X4 FILLER_130_150 ();
 FILLCELL_X4 FILLER_130_158 ();
 FILLCELL_X2 FILLER_130_162 ();
 FILLCELL_X1 FILLER_130_166 ();
 FILLCELL_X2 FILLER_130_205 ();
 FILLCELL_X8 FILLER_130_229 ();
 FILLCELL_X4 FILLER_130_237 ();
 FILLCELL_X1 FILLER_130_262 ();
 FILLCELL_X1 FILLER_130_275 ();
 FILLCELL_X4 FILLER_130_297 ();
 FILLCELL_X1 FILLER_130_301 ();
 FILLCELL_X4 FILLER_130_315 ();
 FILLCELL_X1 FILLER_130_319 ();
 FILLCELL_X4 FILLER_130_378 ();
 FILLCELL_X2 FILLER_130_382 ();
 FILLCELL_X4 FILLER_130_404 ();
 FILLCELL_X2 FILLER_130_408 ();
 FILLCELL_X2 FILLER_130_412 ();
 FILLCELL_X1 FILLER_130_414 ();
 FILLCELL_X8 FILLER_130_423 ();
 FILLCELL_X8 FILLER_130_443 ();
 FILLCELL_X1 FILLER_130_470 ();
 FILLCELL_X2 FILLER_130_475 ();
 FILLCELL_X4 FILLER_130_513 ();
 FILLCELL_X1 FILLER_130_517 ();
 FILLCELL_X8 FILLER_130_552 ();
 FILLCELL_X4 FILLER_130_560 ();
 FILLCELL_X1 FILLER_130_564 ();
 FILLCELL_X2 FILLER_130_569 ();
 FILLCELL_X4 FILLER_130_577 ();
 FILLCELL_X1 FILLER_130_581 ();
 FILLCELL_X4 FILLER_130_584 ();
 FILLCELL_X2 FILLER_130_588 ();
 FILLCELL_X1 FILLER_130_622 ();
 FILLCELL_X1 FILLER_130_626 ();
 FILLCELL_X8 FILLER_130_667 ();
 FILLCELL_X1 FILLER_130_675 ();
 FILLCELL_X2 FILLER_130_679 ();
 FILLCELL_X2 FILLER_130_685 ();
 FILLCELL_X2 FILLER_130_703 ();
 FILLCELL_X1 FILLER_130_707 ();
 FILLCELL_X2 FILLER_130_730 ();
 FILLCELL_X1 FILLER_130_732 ();
 FILLCELL_X1 FILLER_130_735 ();
 FILLCELL_X1 FILLER_130_742 ();
 FILLCELL_X1 FILLER_130_755 ();
 FILLCELL_X1 FILLER_130_760 ();
 FILLCELL_X2 FILLER_130_775 ();
 FILLCELL_X1 FILLER_130_777 ();
 FILLCELL_X4 FILLER_130_798 ();
 FILLCELL_X2 FILLER_130_802 ();
 FILLCELL_X1 FILLER_130_804 ();
 FILLCELL_X4 FILLER_130_815 ();
 FILLCELL_X4 FILLER_130_853 ();
 FILLCELL_X1 FILLER_130_877 ();
 FILLCELL_X1 FILLER_130_898 ();
 FILLCELL_X2 FILLER_130_939 ();
 FILLCELL_X4 FILLER_130_952 ();
 FILLCELL_X1 FILLER_130_956 ();
 FILLCELL_X2 FILLER_130_960 ();
 FILLCELL_X1 FILLER_130_980 ();
 FILLCELL_X1 FILLER_130_987 ();
 FILLCELL_X1 FILLER_130_1003 ();
 FILLCELL_X2 FILLER_130_1011 ();
 FILLCELL_X1 FILLER_130_1013 ();
 FILLCELL_X2 FILLER_130_1017 ();
 FILLCELL_X4 FILLER_130_1054 ();
 FILLCELL_X1 FILLER_130_1068 ();
 FILLCELL_X4 FILLER_130_1094 ();
 FILLCELL_X2 FILLER_130_1098 ();
 FILLCELL_X4 FILLER_131_1 ();
 FILLCELL_X2 FILLER_131_31 ();
 FILLCELL_X4 FILLER_131_37 ();
 FILLCELL_X4 FILLER_131_59 ();
 FILLCELL_X1 FILLER_131_63 ();
 FILLCELL_X1 FILLER_131_82 ();
 FILLCELL_X8 FILLER_131_85 ();
 FILLCELL_X4 FILLER_131_93 ();
 FILLCELL_X1 FILLER_131_97 ();
 FILLCELL_X2 FILLER_131_102 ();
 FILLCELL_X8 FILLER_131_106 ();
 FILLCELL_X4 FILLER_131_114 ();
 FILLCELL_X4 FILLER_131_148 ();
 FILLCELL_X1 FILLER_131_152 ();
 FILLCELL_X8 FILLER_131_173 ();
 FILLCELL_X2 FILLER_131_181 ();
 FILLCELL_X1 FILLER_131_183 ();
 FILLCELL_X8 FILLER_131_186 ();
 FILLCELL_X2 FILLER_131_194 ();
 FILLCELL_X1 FILLER_131_196 ();
 FILLCELL_X8 FILLER_131_219 ();
 FILLCELL_X2 FILLER_131_274 ();
 FILLCELL_X1 FILLER_131_285 ();
 FILLCELL_X4 FILLER_131_290 ();
 FILLCELL_X1 FILLER_131_296 ();
 FILLCELL_X2 FILLER_131_307 ();
 FILLCELL_X2 FILLER_131_313 ();
 FILLCELL_X1 FILLER_131_338 ();
 FILLCELL_X1 FILLER_131_343 ();
 FILLCELL_X4 FILLER_131_366 ();
 FILLCELL_X1 FILLER_131_370 ();
 FILLCELL_X1 FILLER_131_389 ();
 FILLCELL_X2 FILLER_131_392 ();
 FILLCELL_X2 FILLER_131_414 ();
 FILLCELL_X4 FILLER_131_420 ();
 FILLCELL_X2 FILLER_131_424 ();
 FILLCELL_X1 FILLER_131_426 ();
 FILLCELL_X4 FILLER_131_430 ();
 FILLCELL_X2 FILLER_131_434 ();
 FILLCELL_X2 FILLER_131_442 ();
 FILLCELL_X2 FILLER_131_460 ();
 FILLCELL_X1 FILLER_131_464 ();
 FILLCELL_X4 FILLER_131_481 ();
 FILLCELL_X2 FILLER_131_485 ();
 FILLCELL_X8 FILLER_131_491 ();
 FILLCELL_X4 FILLER_131_499 ();
 FILLCELL_X2 FILLER_131_529 ();
 FILLCELL_X1 FILLER_131_531 ();
 FILLCELL_X2 FILLER_131_536 ();
 FILLCELL_X2 FILLER_131_562 ();
 FILLCELL_X1 FILLER_131_564 ();
 FILLCELL_X16 FILLER_131_613 ();
 FILLCELL_X2 FILLER_131_629 ();
 FILLCELL_X1 FILLER_131_637 ();
 FILLCELL_X2 FILLER_131_674 ();
 FILLCELL_X1 FILLER_131_676 ();
 FILLCELL_X2 FILLER_131_681 ();
 FILLCELL_X1 FILLER_131_683 ();
 FILLCELL_X8 FILLER_131_700 ();
 FILLCELL_X1 FILLER_131_708 ();
 FILLCELL_X1 FILLER_131_725 ();
 FILLCELL_X1 FILLER_131_730 ();
 FILLCELL_X1 FILLER_131_741 ();
 FILLCELL_X2 FILLER_131_758 ();
 FILLCELL_X1 FILLER_131_764 ();
 FILLCELL_X8 FILLER_131_769 ();
 FILLCELL_X1 FILLER_131_777 ();
 FILLCELL_X8 FILLER_131_803 ();
 FILLCELL_X2 FILLER_131_811 ();
 FILLCELL_X1 FILLER_131_813 ();
 FILLCELL_X4 FILLER_131_828 ();
 FILLCELL_X4 FILLER_131_835 ();
 FILLCELL_X1 FILLER_131_839 ();
 FILLCELL_X4 FILLER_131_862 ();
 FILLCELL_X1 FILLER_131_866 ();
 FILLCELL_X1 FILLER_131_898 ();
 FILLCELL_X4 FILLER_131_925 ();
 FILLCELL_X2 FILLER_131_929 ();
 FILLCELL_X2 FILLER_131_951 ();
 FILLCELL_X1 FILLER_131_961 ();
 FILLCELL_X1 FILLER_131_997 ();
 FILLCELL_X2 FILLER_131_1016 ();
 FILLCELL_X8 FILLER_131_1032 ();
 FILLCELL_X2 FILLER_131_1040 ();
 FILLCELL_X4 FILLER_131_1098 ();
 FILLCELL_X1 FILLER_131_1102 ();
 FILLCELL_X4 FILLER_132_1 ();
 FILLCELL_X1 FILLER_132_5 ();
 FILLCELL_X2 FILLER_132_14 ();
 FILLCELL_X1 FILLER_132_32 ();
 FILLCELL_X1 FILLER_132_35 ();
 FILLCELL_X1 FILLER_132_104 ();
 FILLCELL_X8 FILLER_132_113 ();
 FILLCELL_X1 FILLER_132_143 ();
 FILLCELL_X4 FILLER_132_164 ();
 FILLCELL_X2 FILLER_132_168 ();
 FILLCELL_X1 FILLER_132_170 ();
 FILLCELL_X16 FILLER_132_205 ();
 FILLCELL_X2 FILLER_132_221 ();
 FILLCELL_X4 FILLER_132_233 ();
 FILLCELL_X1 FILLER_132_237 ();
 FILLCELL_X2 FILLER_132_265 ();
 FILLCELL_X1 FILLER_132_277 ();
 FILLCELL_X4 FILLER_132_305 ();
 FILLCELL_X1 FILLER_132_325 ();
 FILLCELL_X1 FILLER_132_328 ();
 FILLCELL_X8 FILLER_132_345 ();
 FILLCELL_X2 FILLER_132_353 ();
 FILLCELL_X2 FILLER_132_358 ();
 FILLCELL_X1 FILLER_132_360 ();
 FILLCELL_X16 FILLER_132_371 ();
 FILLCELL_X4 FILLER_132_387 ();
 FILLCELL_X2 FILLER_132_391 ();
 FILLCELL_X1 FILLER_132_393 ();
 FILLCELL_X2 FILLER_132_402 ();
 FILLCELL_X1 FILLER_132_404 ();
 FILLCELL_X2 FILLER_132_449 ();
 FILLCELL_X4 FILLER_132_467 ();
 FILLCELL_X2 FILLER_132_471 ();
 FILLCELL_X1 FILLER_132_478 ();
 FILLCELL_X1 FILLER_132_495 ();
 FILLCELL_X1 FILLER_132_500 ();
 FILLCELL_X1 FILLER_132_505 ();
 FILLCELL_X2 FILLER_132_520 ();
 FILLCELL_X2 FILLER_132_546 ();
 FILLCELL_X1 FILLER_132_548 ();
 FILLCELL_X4 FILLER_132_556 ();
 FILLCELL_X2 FILLER_132_560 ();
 FILLCELL_X1 FILLER_132_562 ();
 FILLCELL_X2 FILLER_132_577 ();
 FILLCELL_X2 FILLER_132_583 ();
 FILLCELL_X1 FILLER_132_585 ();
 FILLCELL_X4 FILLER_132_588 ();
 FILLCELL_X1 FILLER_132_592 ();
 FILLCELL_X16 FILLER_132_597 ();
 FILLCELL_X2 FILLER_132_613 ();
 FILLCELL_X1 FILLER_132_668 ();
 FILLCELL_X2 FILLER_132_720 ();
 FILLCELL_X4 FILLER_132_734 ();
 FILLCELL_X2 FILLER_132_738 ();
 FILLCELL_X4 FILLER_132_752 ();
 FILLCELL_X2 FILLER_132_780 ();
 FILLCELL_X8 FILLER_132_802 ();
 FILLCELL_X1 FILLER_132_810 ();
 FILLCELL_X4 FILLER_132_841 ();
 FILLCELL_X2 FILLER_132_845 ();
 FILLCELL_X2 FILLER_132_865 ();
 FILLCELL_X16 FILLER_132_873 ();
 FILLCELL_X4 FILLER_132_916 ();
 FILLCELL_X1 FILLER_132_960 ();
 FILLCELL_X1 FILLER_132_973 ();
 FILLCELL_X4 FILLER_132_981 ();
 FILLCELL_X1 FILLER_132_1001 ();
 FILLCELL_X2 FILLER_132_1055 ();
 FILLCELL_X1 FILLER_132_1059 ();
 FILLCELL_X1 FILLER_132_1070 ();
 FILLCELL_X1 FILLER_132_1127 ();
 FILLCELL_X2 FILLER_133_1 ();
 FILLCELL_X1 FILLER_133_6 ();
 FILLCELL_X8 FILLER_133_13 ();
 FILLCELL_X2 FILLER_133_29 ();
 FILLCELL_X1 FILLER_133_31 ();
 FILLCELL_X2 FILLER_133_46 ();
 FILLCELL_X1 FILLER_133_48 ();
 FILLCELL_X1 FILLER_133_51 ();
 FILLCELL_X1 FILLER_133_56 ();
 FILLCELL_X2 FILLER_133_59 ();
 FILLCELL_X2 FILLER_133_72 ();
 FILLCELL_X1 FILLER_133_74 ();
 FILLCELL_X1 FILLER_133_93 ();
 FILLCELL_X4 FILLER_133_150 ();
 FILLCELL_X1 FILLER_133_164 ();
 FILLCELL_X1 FILLER_133_169 ();
 FILLCELL_X2 FILLER_133_219 ();
 FILLCELL_X1 FILLER_133_221 ();
 FILLCELL_X2 FILLER_133_226 ();
 FILLCELL_X1 FILLER_133_228 ();
 FILLCELL_X2 FILLER_133_233 ();
 FILLCELL_X1 FILLER_133_235 ();
 FILLCELL_X1 FILLER_133_260 ();
 FILLCELL_X4 FILLER_133_271 ();
 FILLCELL_X2 FILLER_133_287 ();
 FILLCELL_X1 FILLER_133_289 ();
 FILLCELL_X2 FILLER_133_303 ();
 FILLCELL_X1 FILLER_133_305 ();
 FILLCELL_X2 FILLER_133_313 ();
 FILLCELL_X1 FILLER_133_363 ();
 FILLCELL_X1 FILLER_133_368 ();
 FILLCELL_X1 FILLER_133_377 ();
 FILLCELL_X2 FILLER_133_416 ();
 FILLCELL_X2 FILLER_133_424 ();
 FILLCELL_X4 FILLER_133_446 ();
 FILLCELL_X2 FILLER_133_450 ();
 FILLCELL_X2 FILLER_133_454 ();
 FILLCELL_X4 FILLER_133_458 ();
 FILLCELL_X2 FILLER_133_508 ();
 FILLCELL_X1 FILLER_133_510 ();
 FILLCELL_X4 FILLER_133_537 ();
 FILLCELL_X2 FILLER_133_541 ();
 FILLCELL_X4 FILLER_133_550 ();
 FILLCELL_X2 FILLER_133_554 ();
 FILLCELL_X1 FILLER_133_556 ();
 FILLCELL_X2 FILLER_133_559 ();
 FILLCELL_X1 FILLER_133_561 ();
 FILLCELL_X1 FILLER_133_586 ();
 FILLCELL_X1 FILLER_133_603 ();
 FILLCELL_X1 FILLER_133_622 ();
 FILLCELL_X8 FILLER_133_625 ();
 FILLCELL_X1 FILLER_133_637 ();
 FILLCELL_X1 FILLER_133_654 ();
 FILLCELL_X1 FILLER_133_663 ();
 FILLCELL_X4 FILLER_133_680 ();
 FILLCELL_X2 FILLER_133_684 ();
 FILLCELL_X1 FILLER_133_686 ();
 FILLCELL_X4 FILLER_133_691 ();
 FILLCELL_X4 FILLER_133_699 ();
 FILLCELL_X2 FILLER_133_703 ();
 FILLCELL_X1 FILLER_133_705 ();
 FILLCELL_X1 FILLER_133_718 ();
 FILLCELL_X2 FILLER_133_763 ();
 FILLCELL_X4 FILLER_133_775 ();
 FILLCELL_X2 FILLER_133_779 ();
 FILLCELL_X1 FILLER_133_801 ();
 FILLCELL_X2 FILLER_133_812 ();
 FILLCELL_X1 FILLER_133_814 ();
 FILLCELL_X2 FILLER_133_831 ();
 FILLCELL_X1 FILLER_133_845 ();
 FILLCELL_X4 FILLER_133_891 ();
 FILLCELL_X1 FILLER_133_906 ();
 FILLCELL_X2 FILLER_133_985 ();
 FILLCELL_X2 FILLER_133_1008 ();
 FILLCELL_X4 FILLER_133_1058 ();
 FILLCELL_X2 FILLER_133_1062 ();
 FILLCELL_X1 FILLER_133_1127 ();
 FILLCELL_X1 FILLER_134_1 ();
 FILLCELL_X1 FILLER_134_18 ();
 FILLCELL_X1 FILLER_134_35 ();
 FILLCELL_X2 FILLER_134_90 ();
 FILLCELL_X2 FILLER_134_110 ();
 FILLCELL_X8 FILLER_134_116 ();
 FILLCELL_X2 FILLER_134_124 ();
 FILLCELL_X1 FILLER_134_146 ();
 FILLCELL_X1 FILLER_134_157 ();
 FILLCELL_X1 FILLER_134_162 ();
 FILLCELL_X2 FILLER_134_173 ();
 FILLCELL_X2 FILLER_134_183 ();
 FILLCELL_X2 FILLER_134_192 ();
 FILLCELL_X1 FILLER_134_289 ();
 FILLCELL_X4 FILLER_134_296 ();
 FILLCELL_X1 FILLER_134_300 ();
 FILLCELL_X2 FILLER_134_312 ();
 FILLCELL_X4 FILLER_134_334 ();
 FILLCELL_X2 FILLER_134_338 ();
 FILLCELL_X2 FILLER_134_342 ();
 FILLCELL_X4 FILLER_134_346 ();
 FILLCELL_X1 FILLER_134_350 ();
 FILLCELL_X4 FILLER_134_381 ();
 FILLCELL_X2 FILLER_134_385 ();
 FILLCELL_X1 FILLER_134_387 ();
 FILLCELL_X2 FILLER_134_391 ();
 FILLCELL_X1 FILLER_134_393 ();
 FILLCELL_X4 FILLER_134_397 ();
 FILLCELL_X2 FILLER_134_401 ();
 FILLCELL_X2 FILLER_134_453 ();
 FILLCELL_X2 FILLER_134_479 ();
 FILLCELL_X1 FILLER_134_487 ();
 FILLCELL_X1 FILLER_134_492 ();
 FILLCELL_X4 FILLER_134_514 ();
 FILLCELL_X1 FILLER_134_518 ();
 FILLCELL_X2 FILLER_134_546 ();
 FILLCELL_X2 FILLER_134_554 ();
 FILLCELL_X1 FILLER_134_556 ();
 FILLCELL_X1 FILLER_134_574 ();
 FILLCELL_X8 FILLER_134_579 ();
 FILLCELL_X4 FILLER_134_587 ();
 FILLCELL_X1 FILLER_134_591 ();
 FILLCELL_X2 FILLER_134_628 ();
 FILLCELL_X1 FILLER_134_630 ();
 FILLCELL_X2 FILLER_134_650 ();
 FILLCELL_X4 FILLER_134_658 ();
 FILLCELL_X2 FILLER_134_665 ();
 FILLCELL_X8 FILLER_134_671 ();
 FILLCELL_X1 FILLER_134_679 ();
 FILLCELL_X4 FILLER_134_682 ();
 FILLCELL_X1 FILLER_134_686 ();
 FILLCELL_X1 FILLER_134_703 ();
 FILLCELL_X1 FILLER_134_728 ();
 FILLCELL_X1 FILLER_134_747 ();
 FILLCELL_X8 FILLER_134_752 ();
 FILLCELL_X4 FILLER_134_760 ();
 FILLCELL_X1 FILLER_134_764 ();
 FILLCELL_X1 FILLER_134_829 ();
 FILLCELL_X1 FILLER_134_846 ();
 FILLCELL_X1 FILLER_134_853 ();
 FILLCELL_X2 FILLER_134_867 ();
 FILLCELL_X8 FILLER_134_893 ();
 FILLCELL_X2 FILLER_134_901 ();
 FILLCELL_X1 FILLER_134_903 ();
 FILLCELL_X1 FILLER_134_911 ();
 FILLCELL_X1 FILLER_134_916 ();
 FILLCELL_X1 FILLER_134_922 ();
 FILLCELL_X1 FILLER_134_928 ();
 FILLCELL_X2 FILLER_134_975 ();
 FILLCELL_X1 FILLER_134_977 ();
 FILLCELL_X1 FILLER_134_985 ();
 FILLCELL_X1 FILLER_134_999 ();
 FILLCELL_X1 FILLER_134_1071 ();
 FILLCELL_X2 FILLER_134_1130 ();
 FILLCELL_X1 FILLER_134_1132 ();
 FILLCELL_X4 FILLER_135_1 ();
 FILLCELL_X2 FILLER_135_5 ();
 FILLCELL_X1 FILLER_135_7 ();
 FILLCELL_X1 FILLER_135_22 ();
 FILLCELL_X1 FILLER_135_27 ();
 FILLCELL_X2 FILLER_135_32 ();
 FILLCELL_X2 FILLER_135_36 ();
 FILLCELL_X1 FILLER_135_38 ();
 FILLCELL_X2 FILLER_135_41 ();
 FILLCELL_X1 FILLER_135_59 ();
 FILLCELL_X2 FILLER_135_76 ();
 FILLCELL_X1 FILLER_135_133 ();
 FILLCELL_X4 FILLER_135_154 ();
 FILLCELL_X1 FILLER_135_178 ();
 FILLCELL_X4 FILLER_135_199 ();
 FILLCELL_X2 FILLER_135_203 ();
 FILLCELL_X1 FILLER_135_205 ();
 FILLCELL_X2 FILLER_135_222 ();
 FILLCELL_X2 FILLER_135_226 ();
 FILLCELL_X4 FILLER_135_257 ();
 FILLCELL_X1 FILLER_135_271 ();
 FILLCELL_X4 FILLER_135_281 ();
 FILLCELL_X4 FILLER_135_298 ();
 FILLCELL_X1 FILLER_135_312 ();
 FILLCELL_X1 FILLER_135_349 ();
 FILLCELL_X2 FILLER_135_398 ();
 FILLCELL_X1 FILLER_135_400 ();
 FILLCELL_X4 FILLER_135_403 ();
 FILLCELL_X1 FILLER_135_411 ();
 FILLCELL_X4 FILLER_135_420 ();
 FILLCELL_X2 FILLER_135_424 ();
 FILLCELL_X2 FILLER_135_432 ();
 FILLCELL_X2 FILLER_135_438 ();
 FILLCELL_X1 FILLER_135_440 ();
 FILLCELL_X2 FILLER_135_445 ();
 FILLCELL_X1 FILLER_135_447 ();
 FILLCELL_X2 FILLER_135_452 ();
 FILLCELL_X4 FILLER_135_470 ();
 FILLCELL_X2 FILLER_135_525 ();
 FILLCELL_X1 FILLER_135_527 ();
 FILLCELL_X2 FILLER_135_551 ();
 FILLCELL_X2 FILLER_135_557 ();
 FILLCELL_X1 FILLER_135_613 ();
 FILLCELL_X1 FILLER_135_630 ();
 FILLCELL_X1 FILLER_135_633 ();
 FILLCELL_X1 FILLER_135_659 ();
 FILLCELL_X1 FILLER_135_700 ();
 FILLCELL_X1 FILLER_135_707 ();
 FILLCELL_X2 FILLER_135_712 ();
 FILLCELL_X2 FILLER_135_718 ();
 FILLCELL_X1 FILLER_135_720 ();
 FILLCELL_X4 FILLER_135_775 ();
 FILLCELL_X1 FILLER_135_779 ();
 FILLCELL_X2 FILLER_135_800 ();
 FILLCELL_X1 FILLER_135_802 ();
 FILLCELL_X1 FILLER_135_806 ();
 FILLCELL_X1 FILLER_135_810 ();
 FILLCELL_X1 FILLER_135_817 ();
 FILLCELL_X2 FILLER_135_830 ();
 FILLCELL_X1 FILLER_135_832 ();
 FILLCELL_X4 FILLER_135_841 ();
 FILLCELL_X16 FILLER_135_869 ();
 FILLCELL_X8 FILLER_135_885 ();
 FILLCELL_X1 FILLER_135_893 ();
 FILLCELL_X4 FILLER_135_898 ();
 FILLCELL_X4 FILLER_135_945 ();
 FILLCELL_X1 FILLER_135_949 ();
 FILLCELL_X1 FILLER_135_990 ();
 FILLCELL_X2 FILLER_135_997 ();
 FILLCELL_X2 FILLER_135_1006 ();
 FILLCELL_X1 FILLER_135_1012 ();
 FILLCELL_X2 FILLER_135_1017 ();
 FILLCELL_X1 FILLER_135_1022 ();
 FILLCELL_X2 FILLER_135_1027 ();
 FILLCELL_X1 FILLER_135_1038 ();
 FILLCELL_X2 FILLER_135_1043 ();
 FILLCELL_X4 FILLER_135_1048 ();
 FILLCELL_X1 FILLER_135_1083 ();
 FILLCELL_X2 FILLER_135_1097 ();
 FILLCELL_X2 FILLER_135_1103 ();
 FILLCELL_X2 FILLER_135_1110 ();
 FILLCELL_X4 FILLER_135_1116 ();
 FILLCELL_X2 FILLER_135_1120 ();
 FILLCELL_X1 FILLER_135_1130 ();
 FILLCELL_X4 FILLER_135_1137 ();
 FILLCELL_X1 FILLER_135_1141 ();
 FILLCELL_X2 FILLER_135_1145 ();
 FILLCELL_X1 FILLER_135_1147 ();
 FILLCELL_X8 FILLER_136_1 ();
 FILLCELL_X1 FILLER_136_9 ();
 FILLCELL_X2 FILLER_136_33 ();
 FILLCELL_X1 FILLER_136_35 ();
 FILLCELL_X1 FILLER_136_40 ();
 FILLCELL_X8 FILLER_136_53 ();
 FILLCELL_X4 FILLER_136_61 ();
 FILLCELL_X8 FILLER_136_83 ();
 FILLCELL_X4 FILLER_136_95 ();
 FILLCELL_X1 FILLER_136_99 ();
 FILLCELL_X8 FILLER_136_116 ();
 FILLCELL_X8 FILLER_136_134 ();
 FILLCELL_X4 FILLER_136_162 ();
 FILLCELL_X2 FILLER_136_166 ();
 FILLCELL_X2 FILLER_136_186 ();
 FILLCELL_X2 FILLER_136_203 ();
 FILLCELL_X1 FILLER_136_205 ();
 FILLCELL_X1 FILLER_136_218 ();
 FILLCELL_X1 FILLER_136_256 ();
 FILLCELL_X1 FILLER_136_261 ();
 FILLCELL_X1 FILLER_136_266 ();
 FILLCELL_X2 FILLER_136_270 ();
 FILLCELL_X2 FILLER_136_275 ();
 FILLCELL_X1 FILLER_136_277 ();
 FILLCELL_X1 FILLER_136_293 ();
 FILLCELL_X1 FILLER_136_298 ();
 FILLCELL_X4 FILLER_136_303 ();
 FILLCELL_X1 FILLER_136_325 ();
 FILLCELL_X2 FILLER_136_330 ();
 FILLCELL_X1 FILLER_136_332 ();
 FILLCELL_X2 FILLER_136_337 ();
 FILLCELL_X1 FILLER_136_339 ();
 FILLCELL_X8 FILLER_136_360 ();
 FILLCELL_X4 FILLER_136_368 ();
 FILLCELL_X2 FILLER_136_372 ();
 FILLCELL_X1 FILLER_136_374 ();
 FILLCELL_X1 FILLER_136_399 ();
 FILLCELL_X1 FILLER_136_410 ();
 FILLCELL_X4 FILLER_136_431 ();
 FILLCELL_X1 FILLER_136_435 ();
 FILLCELL_X1 FILLER_136_438 ();
 FILLCELL_X2 FILLER_136_459 ();
 FILLCELL_X1 FILLER_136_461 ();
 FILLCELL_X1 FILLER_136_480 ();
 FILLCELL_X2 FILLER_136_507 ();
 FILLCELL_X1 FILLER_136_509 ();
 FILLCELL_X1 FILLER_136_512 ();
 FILLCELL_X1 FILLER_136_539 ();
 FILLCELL_X1 FILLER_136_576 ();
 FILLCELL_X2 FILLER_136_579 ();
 FILLCELL_X1 FILLER_136_603 ();
 FILLCELL_X1 FILLER_136_620 ();
 FILLCELL_X1 FILLER_136_625 ();
 FILLCELL_X1 FILLER_136_628 ();
 FILLCELL_X4 FILLER_136_656 ();
 FILLCELL_X8 FILLER_136_702 ();
 FILLCELL_X2 FILLER_136_730 ();
 FILLCELL_X1 FILLER_136_732 ();
 FILLCELL_X4 FILLER_136_747 ();
 FILLCELL_X1 FILLER_136_753 ();
 FILLCELL_X1 FILLER_136_756 ();
 FILLCELL_X2 FILLER_136_761 ();
 FILLCELL_X8 FILLER_136_769 ();
 FILLCELL_X2 FILLER_136_777 ();
 FILLCELL_X1 FILLER_136_779 ();
 FILLCELL_X1 FILLER_136_815 ();
 FILLCELL_X4 FILLER_136_828 ();
 FILLCELL_X2 FILLER_136_832 ();
 FILLCELL_X1 FILLER_136_834 ();
 FILLCELL_X1 FILLER_136_890 ();
 FILLCELL_X1 FILLER_136_905 ();
 FILLCELL_X2 FILLER_136_953 ();
 FILLCELL_X2 FILLER_136_960 ();
 FILLCELL_X1 FILLER_136_979 ();
 FILLCELL_X1 FILLER_136_985 ();
 FILLCELL_X2 FILLER_136_992 ();
 FILLCELL_X1 FILLER_136_1006 ();
 FILLCELL_X1 FILLER_136_1068 ();
 FILLCELL_X2 FILLER_136_1119 ();
 FILLCELL_X1 FILLER_136_1127 ();
 FILLCELL_X1 FILLER_136_1138 ();
 FILLCELL_X16 FILLER_137_1 ();
 FILLCELL_X2 FILLER_137_17 ();
 FILLCELL_X2 FILLER_137_23 ();
 FILLCELL_X2 FILLER_137_29 ();
 FILLCELL_X4 FILLER_137_51 ();
 FILLCELL_X2 FILLER_137_55 ();
 FILLCELL_X1 FILLER_137_57 ();
 FILLCELL_X4 FILLER_137_61 ();
 FILLCELL_X2 FILLER_137_70 ();
 FILLCELL_X1 FILLER_137_72 ();
 FILLCELL_X2 FILLER_137_89 ();
 FILLCELL_X8 FILLER_137_95 ();
 FILLCELL_X4 FILLER_137_103 ();
 FILLCELL_X1 FILLER_137_107 ();
 FILLCELL_X8 FILLER_137_111 ();
 FILLCELL_X8 FILLER_137_141 ();
 FILLCELL_X2 FILLER_137_149 ();
 FILLCELL_X1 FILLER_137_151 ();
 FILLCELL_X1 FILLER_137_160 ();
 FILLCELL_X1 FILLER_137_165 ();
 FILLCELL_X2 FILLER_137_186 ();
 FILLCELL_X8 FILLER_137_230 ();
 FILLCELL_X2 FILLER_137_238 ();
 FILLCELL_X1 FILLER_137_254 ();
 FILLCELL_X4 FILLER_137_268 ();
 FILLCELL_X4 FILLER_137_278 ();
 FILLCELL_X4 FILLER_137_286 ();
 FILLCELL_X1 FILLER_137_290 ();
 FILLCELL_X16 FILLER_137_293 ();
 FILLCELL_X4 FILLER_137_309 ();
 FILLCELL_X1 FILLER_137_313 ();
 FILLCELL_X2 FILLER_137_316 ();
 FILLCELL_X2 FILLER_137_334 ();
 FILLCELL_X4 FILLER_137_354 ();
 FILLCELL_X1 FILLER_137_358 ();
 FILLCELL_X1 FILLER_137_389 ();
 FILLCELL_X1 FILLER_137_392 ();
 FILLCELL_X1 FILLER_137_399 ();
 FILLCELL_X4 FILLER_137_408 ();
 FILLCELL_X2 FILLER_137_412 ();
 FILLCELL_X1 FILLER_137_414 ();
 FILLCELL_X1 FILLER_137_423 ();
 FILLCELL_X1 FILLER_137_466 ();
 FILLCELL_X1 FILLER_137_471 ();
 FILLCELL_X2 FILLER_137_496 ();
 FILLCELL_X1 FILLER_137_498 ();
 FILLCELL_X1 FILLER_137_505 ();
 FILLCELL_X4 FILLER_137_557 ();
 FILLCELL_X2 FILLER_137_565 ();
 FILLCELL_X4 FILLER_137_571 ();
 FILLCELL_X2 FILLER_137_575 ();
 FILLCELL_X4 FILLER_137_579 ();
 FILLCELL_X16 FILLER_137_588 ();
 FILLCELL_X2 FILLER_137_604 ();
 FILLCELL_X1 FILLER_137_606 ();
 FILLCELL_X2 FILLER_137_609 ();
 FILLCELL_X2 FILLER_137_615 ();
 FILLCELL_X1 FILLER_137_649 ();
 FILLCELL_X1 FILLER_137_652 ();
 FILLCELL_X2 FILLER_137_664 ();
 FILLCELL_X1 FILLER_137_669 ();
 FILLCELL_X4 FILLER_137_678 ();
 FILLCELL_X2 FILLER_137_682 ();
 FILLCELL_X1 FILLER_137_684 ();
 FILLCELL_X4 FILLER_137_687 ();
 FILLCELL_X4 FILLER_137_695 ();
 FILLCELL_X1 FILLER_137_699 ();
 FILLCELL_X1 FILLER_137_704 ();
 FILLCELL_X1 FILLER_137_719 ();
 FILLCELL_X2 FILLER_137_725 ();
 FILLCELL_X2 FILLER_137_779 ();
 FILLCELL_X4 FILLER_137_783 ();
 FILLCELL_X2 FILLER_137_787 ();
 FILLCELL_X1 FILLER_137_789 ();
 FILLCELL_X8 FILLER_137_793 ();
 FILLCELL_X2 FILLER_137_801 ();
 FILLCELL_X1 FILLER_137_820 ();
 FILLCELL_X1 FILLER_137_825 ();
 FILLCELL_X2 FILLER_137_848 ();
 FILLCELL_X1 FILLER_137_856 ();
 FILLCELL_X2 FILLER_137_867 ();
 FILLCELL_X1 FILLER_137_869 ();
 FILLCELL_X1 FILLER_137_895 ();
 FILLCELL_X1 FILLER_137_902 ();
 FILLCELL_X1 FILLER_137_910 ();
 FILLCELL_X1 FILLER_137_1106 ();
 FILLCELL_X2 FILLER_137_1117 ();
 FILLCELL_X8 FILLER_137_1138 ();
 FILLCELL_X2 FILLER_137_1146 ();
 FILLCELL_X16 FILLER_138_1 ();
 FILLCELL_X8 FILLER_138_17 ();
 FILLCELL_X2 FILLER_138_35 ();
 FILLCELL_X4 FILLER_138_41 ();
 FILLCELL_X2 FILLER_138_45 ();
 FILLCELL_X2 FILLER_138_49 ();
 FILLCELL_X1 FILLER_138_51 ();
 FILLCELL_X1 FILLER_138_68 ();
 FILLCELL_X1 FILLER_138_71 ();
 FILLCELL_X1 FILLER_138_76 ();
 FILLCELL_X1 FILLER_138_81 ();
 FILLCELL_X2 FILLER_138_104 ();
 FILLCELL_X1 FILLER_138_106 ();
 FILLCELL_X1 FILLER_138_115 ();
 FILLCELL_X1 FILLER_138_138 ();
 FILLCELL_X2 FILLER_138_144 ();
 FILLCELL_X2 FILLER_138_166 ();
 FILLCELL_X2 FILLER_138_213 ();
 FILLCELL_X2 FILLER_138_223 ();
 FILLCELL_X1 FILLER_138_225 ();
 FILLCELL_X2 FILLER_138_247 ();
 FILLCELL_X1 FILLER_138_249 ();
 FILLCELL_X1 FILLER_138_253 ();
 FILLCELL_X32 FILLER_138_276 ();
 FILLCELL_X16 FILLER_138_308 ();
 FILLCELL_X8 FILLER_138_324 ();
 FILLCELL_X4 FILLER_138_332 ();
 FILLCELL_X4 FILLER_138_352 ();
 FILLCELL_X8 FILLER_138_380 ();
 FILLCELL_X2 FILLER_138_477 ();
 FILLCELL_X4 FILLER_138_550 ();
 FILLCELL_X1 FILLER_138_554 ();
 FILLCELL_X2 FILLER_138_558 ();
 FILLCELL_X2 FILLER_138_576 ();
 FILLCELL_X2 FILLER_138_594 ();
 FILLCELL_X2 FILLER_138_602 ();
 FILLCELL_X1 FILLER_138_604 ();
 FILLCELL_X1 FILLER_138_621 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X2 FILLER_138_632 ();
 FILLCELL_X1 FILLER_138_634 ();
 FILLCELL_X2 FILLER_138_653 ();
 FILLCELL_X2 FILLER_138_657 ();
 FILLCELL_X4 FILLER_138_686 ();
 FILLCELL_X1 FILLER_138_715 ();
 FILLCELL_X4 FILLER_138_736 ();
 FILLCELL_X2 FILLER_138_740 ();
 FILLCELL_X1 FILLER_138_742 ();
 FILLCELL_X1 FILLER_138_745 ();
 FILLCELL_X2 FILLER_138_766 ();
 FILLCELL_X1 FILLER_138_808 ();
 FILLCELL_X2 FILLER_138_824 ();
 FILLCELL_X4 FILLER_138_832 ();
 FILLCELL_X2 FILLER_138_836 ();
 FILLCELL_X1 FILLER_138_840 ();
 FILLCELL_X2 FILLER_138_868 ();
 FILLCELL_X1 FILLER_138_913 ();
 FILLCELL_X1 FILLER_138_924 ();
 FILLCELL_X1 FILLER_138_929 ();
 FILLCELL_X2 FILLER_138_966 ();
 FILLCELL_X1 FILLER_138_968 ();
 FILLCELL_X1 FILLER_138_1017 ();
 FILLCELL_X1 FILLER_138_1066 ();
 FILLCELL_X1 FILLER_138_1078 ();
 FILLCELL_X1 FILLER_138_1090 ();
 FILLCELL_X1 FILLER_138_1096 ();
 FILLCELL_X1 FILLER_138_1104 ();
 FILLCELL_X1 FILLER_138_1123 ();
 FILLCELL_X1 FILLER_138_1128 ();
 FILLCELL_X1 FILLER_138_1136 ();
 FILLCELL_X1 FILLER_138_1147 ();
 FILLCELL_X16 FILLER_139_1 ();
 FILLCELL_X8 FILLER_139_17 ();
 FILLCELL_X2 FILLER_139_25 ();
 FILLCELL_X4 FILLER_139_31 ();
 FILLCELL_X2 FILLER_139_35 ();
 FILLCELL_X4 FILLER_139_41 ();
 FILLCELL_X2 FILLER_139_67 ();
 FILLCELL_X4 FILLER_139_85 ();
 FILLCELL_X1 FILLER_139_97 ();
 FILLCELL_X8 FILLER_139_100 ();
 FILLCELL_X1 FILLER_139_108 ();
 FILLCELL_X2 FILLER_139_129 ();
 FILLCELL_X8 FILLER_139_150 ();
 FILLCELL_X1 FILLER_139_158 ();
 FILLCELL_X1 FILLER_139_163 ();
 FILLCELL_X1 FILLER_139_168 ();
 FILLCELL_X1 FILLER_139_173 ();
 FILLCELL_X4 FILLER_139_184 ();
 FILLCELL_X1 FILLER_139_188 ();
 FILLCELL_X1 FILLER_139_233 ();
 FILLCELL_X1 FILLER_139_238 ();
 FILLCELL_X1 FILLER_139_246 ();
 FILLCELL_X2 FILLER_139_251 ();
 FILLCELL_X1 FILLER_139_263 ();
 FILLCELL_X32 FILLER_139_271 ();
 FILLCELL_X4 FILLER_139_303 ();
 FILLCELL_X2 FILLER_139_307 ();
 FILLCELL_X8 FILLER_139_329 ();
 FILLCELL_X2 FILLER_139_337 ();
 FILLCELL_X1 FILLER_139_339 ();
 FILLCELL_X4 FILLER_139_356 ();
 FILLCELL_X2 FILLER_139_360 ();
 FILLCELL_X1 FILLER_139_362 ();
 FILLCELL_X4 FILLER_139_369 ();
 FILLCELL_X1 FILLER_139_373 ();
 FILLCELL_X2 FILLER_139_402 ();
 FILLCELL_X2 FILLER_139_461 ();
 FILLCELL_X1 FILLER_139_463 ();
 FILLCELL_X2 FILLER_139_478 ();
 FILLCELL_X1 FILLER_139_484 ();
 FILLCELL_X2 FILLER_139_523 ();
 FILLCELL_X1 FILLER_139_529 ();
 FILLCELL_X2 FILLER_139_565 ();
 FILLCELL_X2 FILLER_139_571 ();
 FILLCELL_X2 FILLER_139_577 ();
 FILLCELL_X2 FILLER_139_583 ();
 FILLCELL_X2 FILLER_139_589 ();
 FILLCELL_X1 FILLER_139_591 ();
 FILLCELL_X4 FILLER_139_606 ();
 FILLCELL_X2 FILLER_139_610 ();
 FILLCELL_X1 FILLER_139_612 ();
 FILLCELL_X4 FILLER_139_615 ();
 FILLCELL_X1 FILLER_139_621 ();
 FILLCELL_X2 FILLER_139_624 ();
 FILLCELL_X1 FILLER_139_626 ();
 FILLCELL_X8 FILLER_139_629 ();
 FILLCELL_X4 FILLER_139_637 ();
 FILLCELL_X2 FILLER_139_641 ();
 FILLCELL_X1 FILLER_139_643 ();
 FILLCELL_X2 FILLER_139_648 ();
 FILLCELL_X4 FILLER_139_664 ();
 FILLCELL_X1 FILLER_139_668 ();
 FILLCELL_X2 FILLER_139_673 ();
 FILLCELL_X1 FILLER_139_675 ();
 FILLCELL_X4 FILLER_139_682 ();
 FILLCELL_X2 FILLER_139_686 ();
 FILLCELL_X4 FILLER_139_692 ();
 FILLCELL_X2 FILLER_139_696 ();
 FILLCELL_X1 FILLER_139_698 ();
 FILLCELL_X1 FILLER_139_706 ();
 FILLCELL_X8 FILLER_139_727 ();
 FILLCELL_X1 FILLER_139_735 ();
 FILLCELL_X8 FILLER_139_738 ();
 FILLCELL_X1 FILLER_139_746 ();
 FILLCELL_X1 FILLER_139_749 ();
 FILLCELL_X4 FILLER_139_770 ();
 FILLCELL_X1 FILLER_139_813 ();
 FILLCELL_X1 FILLER_139_816 ();
 FILLCELL_X1 FILLER_139_825 ();
 FILLCELL_X2 FILLER_139_831 ();
 FILLCELL_X1 FILLER_139_843 ();
 FILLCELL_X1 FILLER_139_858 ();
 FILLCELL_X2 FILLER_139_907 ();
 FILLCELL_X1 FILLER_139_961 ();
 FILLCELL_X1 FILLER_139_965 ();
 FILLCELL_X1 FILLER_139_969 ();
 FILLCELL_X2 FILLER_139_979 ();
 FILLCELL_X2 FILLER_139_1007 ();
 FILLCELL_X1 FILLER_139_1049 ();
 FILLCELL_X1 FILLER_139_1088 ();
 FILLCELL_X2 FILLER_139_1128 ();
 FILLCELL_X4 FILLER_139_1137 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X4 FILLER_140_49 ();
 FILLCELL_X2 FILLER_140_71 ();
 FILLCELL_X1 FILLER_140_73 ();
 FILLCELL_X1 FILLER_140_78 ();
 FILLCELL_X1 FILLER_140_83 ();
 FILLCELL_X4 FILLER_140_100 ();
 FILLCELL_X1 FILLER_140_104 ();
 FILLCELL_X2 FILLER_140_119 ();
 FILLCELL_X1 FILLER_140_137 ();
 FILLCELL_X4 FILLER_140_173 ();
 FILLCELL_X2 FILLER_140_179 ();
 FILLCELL_X8 FILLER_140_183 ();
 FILLCELL_X2 FILLER_140_191 ();
 FILLCELL_X1 FILLER_140_193 ();
 FILLCELL_X1 FILLER_140_217 ();
 FILLCELL_X32 FILLER_140_277 ();
 FILLCELL_X8 FILLER_140_309 ();
 FILLCELL_X1 FILLER_140_317 ();
 FILLCELL_X1 FILLER_140_320 ();
 FILLCELL_X8 FILLER_140_341 ();
 FILLCELL_X1 FILLER_140_349 ();
 FILLCELL_X1 FILLER_140_380 ();
 FILLCELL_X8 FILLER_140_383 ();
 FILLCELL_X1 FILLER_140_391 ();
 FILLCELL_X2 FILLER_140_456 ();
 FILLCELL_X1 FILLER_140_458 ();
 FILLCELL_X8 FILLER_140_463 ();
 FILLCELL_X1 FILLER_140_481 ();
 FILLCELL_X4 FILLER_140_519 ();
 FILLCELL_X1 FILLER_140_530 ();
 FILLCELL_X1 FILLER_140_546 ();
 FILLCELL_X1 FILLER_140_554 ();
 FILLCELL_X2 FILLER_140_560 ();
 FILLCELL_X2 FILLER_140_568 ();
 FILLCELL_X1 FILLER_140_570 ();
 FILLCELL_X2 FILLER_140_574 ();
 FILLCELL_X1 FILLER_140_580 ();
 FILLCELL_X1 FILLER_140_597 ();
 FILLCELL_X1 FILLER_140_614 ();
 FILLCELL_X1 FILLER_140_632 ();
 FILLCELL_X1 FILLER_140_639 ();
 FILLCELL_X4 FILLER_140_658 ();
 FILLCELL_X1 FILLER_140_662 ();
 FILLCELL_X1 FILLER_140_679 ();
 FILLCELL_X1 FILLER_140_700 ();
 FILLCELL_X2 FILLER_140_705 ();
 FILLCELL_X8 FILLER_140_711 ();
 FILLCELL_X2 FILLER_140_727 ();
 FILLCELL_X1 FILLER_140_729 ();
 FILLCELL_X2 FILLER_140_746 ();
 FILLCELL_X8 FILLER_140_750 ();
 FILLCELL_X4 FILLER_140_758 ();
 FILLCELL_X2 FILLER_140_762 ();
 FILLCELL_X1 FILLER_140_784 ();
 FILLCELL_X1 FILLER_140_799 ();
 FILLCELL_X2 FILLER_140_806 ();
 FILLCELL_X1 FILLER_140_808 ();
 FILLCELL_X4 FILLER_140_815 ();
 FILLCELL_X1 FILLER_140_822 ();
 FILLCELL_X1 FILLER_140_827 ();
 FILLCELL_X1 FILLER_140_832 ();
 FILLCELL_X4 FILLER_140_839 ();
 FILLCELL_X1 FILLER_140_849 ();
 FILLCELL_X1 FILLER_140_865 ();
 FILLCELL_X1 FILLER_140_869 ();
 FILLCELL_X1 FILLER_140_873 ();
 FILLCELL_X1 FILLER_140_877 ();
 FILLCELL_X2 FILLER_140_885 ();
 FILLCELL_X1 FILLER_140_907 ();
 FILLCELL_X4 FILLER_140_912 ();
 FILLCELL_X1 FILLER_140_926 ();
 FILLCELL_X1 FILLER_140_1007 ();
 FILLCELL_X1 FILLER_140_1012 ();
 FILLCELL_X2 FILLER_140_1029 ();
 FILLCELL_X1 FILLER_140_1039 ();
 FILLCELL_X2 FILLER_140_1047 ();
 FILLCELL_X1 FILLER_140_1114 ();
 FILLCELL_X16 FILLER_140_1130 ();
 FILLCELL_X2 FILLER_140_1146 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X16 FILLER_141_33 ();
 FILLCELL_X4 FILLER_141_51 ();
 FILLCELL_X2 FILLER_141_55 ();
 FILLCELL_X1 FILLER_141_57 ();
 FILLCELL_X1 FILLER_141_62 ();
 FILLCELL_X4 FILLER_141_69 ();
 FILLCELL_X2 FILLER_141_77 ();
 FILLCELL_X2 FILLER_141_93 ();
 FILLCELL_X1 FILLER_141_95 ();
 FILLCELL_X8 FILLER_141_98 ();
 FILLCELL_X1 FILLER_141_106 ();
 FILLCELL_X1 FILLER_141_111 ();
 FILLCELL_X1 FILLER_141_114 ();
 FILLCELL_X1 FILLER_141_117 ();
 FILLCELL_X1 FILLER_141_122 ();
 FILLCELL_X2 FILLER_141_139 ();
 FILLCELL_X2 FILLER_141_149 ();
 FILLCELL_X2 FILLER_141_155 ();
 FILLCELL_X4 FILLER_141_167 ();
 FILLCELL_X1 FILLER_141_171 ();
 FILLCELL_X1 FILLER_141_190 ();
 FILLCELL_X2 FILLER_141_193 ();
 FILLCELL_X1 FILLER_141_197 ();
 FILLCELL_X1 FILLER_141_228 ();
 FILLCELL_X1 FILLER_141_232 ();
 FILLCELL_X1 FILLER_141_258 ();
 FILLCELL_X1 FILLER_141_262 ();
 FILLCELL_X4 FILLER_141_273 ();
 FILLCELL_X2 FILLER_141_277 ();
 FILLCELL_X16 FILLER_141_283 ();
 FILLCELL_X8 FILLER_141_299 ();
 FILLCELL_X4 FILLER_141_307 ();
 FILLCELL_X4 FILLER_141_313 ();
 FILLCELL_X4 FILLER_141_337 ();
 FILLCELL_X2 FILLER_141_341 ();
 FILLCELL_X16 FILLER_141_389 ();
 FILLCELL_X2 FILLER_141_405 ();
 FILLCELL_X1 FILLER_141_407 ();
 FILLCELL_X2 FILLER_141_410 ();
 FILLCELL_X1 FILLER_141_412 ();
 FILLCELL_X8 FILLER_141_435 ();
 FILLCELL_X4 FILLER_141_463 ();
 FILLCELL_X1 FILLER_141_467 ();
 FILLCELL_X1 FILLER_141_478 ();
 FILLCELL_X1 FILLER_141_489 ();
 FILLCELL_X1 FILLER_141_522 ();
 FILLCELL_X2 FILLER_141_530 ();
 FILLCELL_X2 FILLER_141_535 ();
 FILLCELL_X2 FILLER_141_559 ();
 FILLCELL_X1 FILLER_141_561 ();
 FILLCELL_X2 FILLER_141_568 ();
 FILLCELL_X1 FILLER_141_570 ();
 FILLCELL_X1 FILLER_141_577 ();
 FILLCELL_X2 FILLER_141_587 ();
 FILLCELL_X1 FILLER_141_601 ();
 FILLCELL_X1 FILLER_141_606 ();
 FILLCELL_X1 FILLER_141_623 ();
 FILLCELL_X1 FILLER_141_628 ();
 FILLCELL_X2 FILLER_141_649 ();
 FILLCELL_X2 FILLER_141_659 ();
 FILLCELL_X1 FILLER_141_661 ();
 FILLCELL_X2 FILLER_141_670 ();
 FILLCELL_X1 FILLER_141_672 ();
 FILLCELL_X2 FILLER_141_677 ();
 FILLCELL_X1 FILLER_141_679 ();
 FILLCELL_X2 FILLER_141_694 ();
 FILLCELL_X1 FILLER_141_708 ();
 FILLCELL_X4 FILLER_141_737 ();
 FILLCELL_X1 FILLER_141_741 ();
 FILLCELL_X16 FILLER_141_744 ();
 FILLCELL_X4 FILLER_141_794 ();
 FILLCELL_X2 FILLER_141_832 ();
 FILLCELL_X1 FILLER_141_840 ();
 FILLCELL_X2 FILLER_141_853 ();
 FILLCELL_X4 FILLER_141_867 ();
 FILLCELL_X2 FILLER_141_878 ();
 FILLCELL_X4 FILLER_141_883 ();
 FILLCELL_X1 FILLER_141_887 ();
 FILLCELL_X1 FILLER_141_908 ();
 FILLCELL_X1 FILLER_141_916 ();
 FILLCELL_X1 FILLER_141_924 ();
 FILLCELL_X1 FILLER_141_929 ();
 FILLCELL_X1 FILLER_141_934 ();
 FILLCELL_X4 FILLER_141_944 ();
 FILLCELL_X2 FILLER_141_948 ();
 FILLCELL_X1 FILLER_141_950 ();
 FILLCELL_X2 FILLER_141_956 ();
 FILLCELL_X1 FILLER_141_958 ();
 FILLCELL_X2 FILLER_141_981 ();
 FILLCELL_X1 FILLER_141_1040 ();
 FILLCELL_X1 FILLER_141_1044 ();
 FILLCELL_X2 FILLER_141_1076 ();
 FILLCELL_X1 FILLER_141_1078 ();
 FILLCELL_X2 FILLER_141_1122 ();
 FILLCELL_X16 FILLER_141_1131 ();
 FILLCELL_X1 FILLER_141_1147 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X16 FILLER_142_33 ();
 FILLCELL_X4 FILLER_142_49 ();
 FILLCELL_X2 FILLER_142_53 ();
 FILLCELL_X1 FILLER_142_55 ();
 FILLCELL_X1 FILLER_142_120 ();
 FILLCELL_X1 FILLER_142_123 ();
 FILLCELL_X8 FILLER_142_126 ();
 FILLCELL_X2 FILLER_142_134 ();
 FILLCELL_X2 FILLER_142_172 ();
 FILLCELL_X4 FILLER_142_176 ();
 FILLCELL_X2 FILLER_142_180 ();
 FILLCELL_X1 FILLER_142_182 ();
 FILLCELL_X2 FILLER_142_199 ();
 FILLCELL_X1 FILLER_142_201 ();
 FILLCELL_X16 FILLER_142_204 ();
 FILLCELL_X8 FILLER_142_224 ();
 FILLCELL_X2 FILLER_142_232 ();
 FILLCELL_X1 FILLER_142_234 ();
 FILLCELL_X4 FILLER_142_265 ();
 FILLCELL_X1 FILLER_142_269 ();
 FILLCELL_X16 FILLER_142_294 ();
 FILLCELL_X8 FILLER_142_310 ();
 FILLCELL_X2 FILLER_142_318 ();
 FILLCELL_X4 FILLER_142_322 ();
 FILLCELL_X1 FILLER_142_326 ();
 FILLCELL_X4 FILLER_142_329 ();
 FILLCELL_X2 FILLER_142_333 ();
 FILLCELL_X1 FILLER_142_356 ();
 FILLCELL_X8 FILLER_142_377 ();
 FILLCELL_X4 FILLER_142_385 ();
 FILLCELL_X1 FILLER_142_389 ();
 FILLCELL_X4 FILLER_142_394 ();
 FILLCELL_X2 FILLER_142_398 ();
 FILLCELL_X2 FILLER_142_436 ();
 FILLCELL_X4 FILLER_142_440 ();
 FILLCELL_X2 FILLER_142_494 ();
 FILLCELL_X1 FILLER_142_498 ();
 FILLCELL_X2 FILLER_142_515 ();
 FILLCELL_X1 FILLER_142_517 ();
 FILLCELL_X2 FILLER_142_541 ();
 FILLCELL_X1 FILLER_142_547 ();
 FILLCELL_X2 FILLER_142_590 ();
 FILLCELL_X2 FILLER_142_594 ();
 FILLCELL_X1 FILLER_142_596 ();
 FILLCELL_X2 FILLER_142_616 ();
 FILLCELL_X2 FILLER_142_622 ();
 FILLCELL_X4 FILLER_142_627 ();
 FILLCELL_X4 FILLER_142_635 ();
 FILLCELL_X4 FILLER_142_642 ();
 FILLCELL_X4 FILLER_142_722 ();
 FILLCELL_X1 FILLER_142_726 ();
 FILLCELL_X4 FILLER_142_745 ();
 FILLCELL_X4 FILLER_142_751 ();
 FILLCELL_X1 FILLER_142_755 ();
 FILLCELL_X16 FILLER_142_778 ();
 FILLCELL_X1 FILLER_142_794 ();
 FILLCELL_X2 FILLER_142_817 ();
 FILLCELL_X1 FILLER_142_819 ();
 FILLCELL_X1 FILLER_142_841 ();
 FILLCELL_X1 FILLER_142_847 ();
 FILLCELL_X4 FILLER_142_852 ();
 FILLCELL_X1 FILLER_142_861 ();
 FILLCELL_X1 FILLER_142_868 ();
 FILLCELL_X1 FILLER_142_875 ();
 FILLCELL_X1 FILLER_142_881 ();
 FILLCELL_X16 FILLER_142_887 ();
 FILLCELL_X4 FILLER_142_903 ();
 FILLCELL_X1 FILLER_142_907 ();
 FILLCELL_X1 FILLER_142_928 ();
 FILLCELL_X1 FILLER_142_932 ();
 FILLCELL_X1 FILLER_142_947 ();
 FILLCELL_X1 FILLER_142_957 ();
 FILLCELL_X1 FILLER_142_988 ();
 FILLCELL_X1 FILLER_142_992 ();
 FILLCELL_X1 FILLER_142_999 ();
 FILLCELL_X1 FILLER_142_1009 ();
 FILLCELL_X2 FILLER_142_1047 ();
 FILLCELL_X2 FILLER_142_1098 ();
 FILLCELL_X1 FILLER_142_1100 ();
 FILLCELL_X16 FILLER_142_1120 ();
 FILLCELL_X8 FILLER_142_1136 ();
 FILLCELL_X4 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X16 FILLER_143_33 ();
 FILLCELL_X8 FILLER_143_49 ();
 FILLCELL_X1 FILLER_143_57 ();
 FILLCELL_X8 FILLER_143_76 ();
 FILLCELL_X1 FILLER_143_84 ();
 FILLCELL_X4 FILLER_143_105 ();
 FILLCELL_X2 FILLER_143_109 ();
 FILLCELL_X1 FILLER_143_111 ();
 FILLCELL_X2 FILLER_143_131 ();
 FILLCELL_X2 FILLER_143_149 ();
 FILLCELL_X2 FILLER_143_153 ();
 FILLCELL_X1 FILLER_143_155 ();
 FILLCELL_X8 FILLER_143_158 ();
 FILLCELL_X1 FILLER_143_166 ();
 FILLCELL_X16 FILLER_143_183 ();
 FILLCELL_X4 FILLER_143_199 ();
 FILLCELL_X4 FILLER_143_233 ();
 FILLCELL_X2 FILLER_143_237 ();
 FILLCELL_X32 FILLER_143_259 ();
 FILLCELL_X16 FILLER_143_291 ();
 FILLCELL_X1 FILLER_143_307 ();
 FILLCELL_X1 FILLER_143_391 ();
 FILLCELL_X8 FILLER_143_431 ();
 FILLCELL_X4 FILLER_143_439 ();
 FILLCELL_X2 FILLER_143_443 ();
 FILLCELL_X16 FILLER_143_447 ();
 FILLCELL_X1 FILLER_143_463 ();
 FILLCELL_X2 FILLER_143_466 ();
 FILLCELL_X1 FILLER_143_535 ();
 FILLCELL_X2 FILLER_143_577 ();
 FILLCELL_X1 FILLER_143_579 ();
 FILLCELL_X1 FILLER_143_603 ();
 FILLCELL_X2 FILLER_143_607 ();
 FILLCELL_X2 FILLER_143_668 ();
 FILLCELL_X2 FILLER_143_678 ();
 FILLCELL_X1 FILLER_143_680 ();
 FILLCELL_X4 FILLER_143_700 ();
 FILLCELL_X4 FILLER_143_706 ();
 FILLCELL_X2 FILLER_143_710 ();
 FILLCELL_X2 FILLER_143_724 ();
 FILLCELL_X2 FILLER_143_796 ();
 FILLCELL_X1 FILLER_143_833 ();
 FILLCELL_X8 FILLER_143_836 ();
 FILLCELL_X4 FILLER_143_844 ();
 FILLCELL_X1 FILLER_143_848 ();
 FILLCELL_X4 FILLER_143_855 ();
 FILLCELL_X2 FILLER_143_859 ();
 FILLCELL_X8 FILLER_143_865 ();
 FILLCELL_X2 FILLER_143_873 ();
 FILLCELL_X32 FILLER_143_889 ();
 FILLCELL_X4 FILLER_143_921 ();
 FILLCELL_X2 FILLER_143_945 ();
 FILLCELL_X2 FILLER_143_1000 ();
 FILLCELL_X1 FILLER_143_1015 ();
 FILLCELL_X1 FILLER_143_1031 ();
 FILLCELL_X1 FILLER_143_1098 ();
 FILLCELL_X16 FILLER_143_1122 ();
 FILLCELL_X8 FILLER_143_1138 ();
 FILLCELL_X2 FILLER_143_1146 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X8 FILLER_144_65 ();
 FILLCELL_X2 FILLER_144_73 ();
 FILLCELL_X8 FILLER_144_95 ();
 FILLCELL_X2 FILLER_144_103 ();
 FILLCELL_X8 FILLER_144_142 ();
 FILLCELL_X8 FILLER_144_166 ();
 FILLCELL_X1 FILLER_144_174 ();
 FILLCELL_X4 FILLER_144_177 ();
 FILLCELL_X4 FILLER_144_185 ();
 FILLCELL_X2 FILLER_144_189 ();
 FILLCELL_X1 FILLER_144_191 ();
 FILLCELL_X4 FILLER_144_216 ();
 FILLCELL_X32 FILLER_144_258 ();
 FILLCELL_X8 FILLER_144_290 ();
 FILLCELL_X4 FILLER_144_298 ();
 FILLCELL_X2 FILLER_144_302 ();
 FILLCELL_X4 FILLER_144_322 ();
 FILLCELL_X1 FILLER_144_326 ();
 FILLCELL_X1 FILLER_144_334 ();
 FILLCELL_X2 FILLER_144_340 ();
 FILLCELL_X2 FILLER_144_364 ();
 FILLCELL_X1 FILLER_144_366 ();
 FILLCELL_X1 FILLER_144_402 ();
 FILLCELL_X2 FILLER_144_437 ();
 FILLCELL_X8 FILLER_144_455 ();
 FILLCELL_X2 FILLER_144_463 ();
 FILLCELL_X4 FILLER_144_487 ();
 FILLCELL_X2 FILLER_144_491 ();
 FILLCELL_X1 FILLER_144_493 ();
 FILLCELL_X1 FILLER_144_553 ();
 FILLCELL_X8 FILLER_144_564 ();
 FILLCELL_X1 FILLER_144_576 ();
 FILLCELL_X1 FILLER_144_581 ();
 FILLCELL_X1 FILLER_144_588 ();
 FILLCELL_X1 FILLER_144_609 ();
 FILLCELL_X2 FILLER_144_613 ();
 FILLCELL_X1 FILLER_144_615 ();
 FILLCELL_X1 FILLER_144_619 ();
 FILLCELL_X4 FILLER_144_626 ();
 FILLCELL_X1 FILLER_144_630 ();
 FILLCELL_X8 FILLER_144_632 ();
 FILLCELL_X2 FILLER_144_640 ();
 FILLCELL_X1 FILLER_144_642 ();
 FILLCELL_X4 FILLER_144_645 ();
 FILLCELL_X1 FILLER_144_649 ();
 FILLCELL_X2 FILLER_144_654 ();
 FILLCELL_X4 FILLER_144_658 ();
 FILLCELL_X8 FILLER_144_682 ();
 FILLCELL_X4 FILLER_144_690 ();
 FILLCELL_X2 FILLER_144_694 ();
 FILLCELL_X1 FILLER_144_696 ();
 FILLCELL_X4 FILLER_144_706 ();
 FILLCELL_X8 FILLER_144_730 ();
 FILLCELL_X4 FILLER_144_738 ();
 FILLCELL_X2 FILLER_144_742 ();
 FILLCELL_X1 FILLER_144_744 ();
 FILLCELL_X2 FILLER_144_763 ();
 FILLCELL_X2 FILLER_144_785 ();
 FILLCELL_X1 FILLER_144_787 ();
 FILLCELL_X2 FILLER_144_802 ();
 FILLCELL_X2 FILLER_144_806 ();
 FILLCELL_X1 FILLER_144_808 ();
 FILLCELL_X1 FILLER_144_882 ();
 FILLCELL_X16 FILLER_144_893 ();
 FILLCELL_X8 FILLER_144_909 ();
 FILLCELL_X4 FILLER_144_917 ();
 FILLCELL_X4 FILLER_144_941 ();
 FILLCELL_X1 FILLER_144_945 ();
 FILLCELL_X2 FILLER_144_952 ();
 FILLCELL_X1 FILLER_144_961 ();
 FILLCELL_X4 FILLER_144_975 ();
 FILLCELL_X1 FILLER_144_979 ();
 FILLCELL_X1 FILLER_144_991 ();
 FILLCELL_X1 FILLER_144_996 ();
 FILLCELL_X1 FILLER_144_1004 ();
 FILLCELL_X1 FILLER_144_1011 ();
 FILLCELL_X2 FILLER_144_1098 ();
 FILLCELL_X32 FILLER_144_1110 ();
 FILLCELL_X4 FILLER_144_1142 ();
 FILLCELL_X2 FILLER_144_1146 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X4 FILLER_145_65 ();
 FILLCELL_X1 FILLER_145_69 ();
 FILLCELL_X8 FILLER_145_112 ();
 FILLCELL_X2 FILLER_145_122 ();
 FILLCELL_X4 FILLER_145_134 ();
 FILLCELL_X1 FILLER_145_138 ();
 FILLCELL_X2 FILLER_145_141 ();
 FILLCELL_X32 FILLER_145_250 ();
 FILLCELL_X32 FILLER_145_282 ();
 FILLCELL_X4 FILLER_145_314 ();
 FILLCELL_X2 FILLER_145_318 ();
 FILLCELL_X4 FILLER_145_338 ();
 FILLCELL_X2 FILLER_145_342 ();
 FILLCELL_X1 FILLER_145_344 ();
 FILLCELL_X2 FILLER_145_347 ();
 FILLCELL_X1 FILLER_145_349 ();
 FILLCELL_X4 FILLER_145_353 ();
 FILLCELL_X1 FILLER_145_357 ();
 FILLCELL_X2 FILLER_145_378 ();
 FILLCELL_X16 FILLER_145_382 ();
 FILLCELL_X8 FILLER_145_398 ();
 FILLCELL_X4 FILLER_145_406 ();
 FILLCELL_X2 FILLER_145_410 ();
 FILLCELL_X1 FILLER_145_414 ();
 FILLCELL_X1 FILLER_145_417 ();
 FILLCELL_X1 FILLER_145_425 ();
 FILLCELL_X1 FILLER_145_442 ();
 FILLCELL_X8 FILLER_145_447 ();
 FILLCELL_X2 FILLER_145_455 ();
 FILLCELL_X1 FILLER_145_457 ();
 FILLCELL_X2 FILLER_145_474 ();
 FILLCELL_X4 FILLER_145_498 ();
 FILLCELL_X1 FILLER_145_502 ();
 FILLCELL_X1 FILLER_145_568 ();
 FILLCELL_X2 FILLER_145_579 ();
 FILLCELL_X1 FILLER_145_601 ();
 FILLCELL_X1 FILLER_145_647 ();
 FILLCELL_X2 FILLER_145_664 ();
 FILLCELL_X1 FILLER_145_666 ();
 FILLCELL_X4 FILLER_145_670 ();
 FILLCELL_X2 FILLER_145_756 ();
 FILLCELL_X1 FILLER_145_758 ();
 FILLCELL_X1 FILLER_145_768 ();
 FILLCELL_X8 FILLER_145_789 ();
 FILLCELL_X2 FILLER_145_797 ();
 FILLCELL_X1 FILLER_145_799 ();
 FILLCELL_X2 FILLER_145_806 ();
 FILLCELL_X1 FILLER_145_808 ();
 FILLCELL_X1 FILLER_145_882 ();
 FILLCELL_X32 FILLER_145_887 ();
 FILLCELL_X32 FILLER_145_919 ();
 FILLCELL_X2 FILLER_145_951 ();
 FILLCELL_X2 FILLER_145_964 ();
 FILLCELL_X4 FILLER_145_974 ();
 FILLCELL_X1 FILLER_145_1009 ();
 FILLCELL_X1 FILLER_145_1020 ();
 FILLCELL_X2 FILLER_145_1034 ();
 FILLCELL_X1 FILLER_145_1053 ();
 FILLCELL_X1 FILLER_145_1064 ();
 FILLCELL_X1 FILLER_145_1094 ();
 FILLCELL_X4 FILLER_145_1098 ();
 FILLCELL_X32 FILLER_145_1109 ();
 FILLCELL_X4 FILLER_145_1141 ();
 FILLCELL_X2 FILLER_145_1145 ();
 FILLCELL_X1 FILLER_145_1147 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X8 FILLER_146_97 ();
 FILLCELL_X2 FILLER_146_105 ();
 FILLCELL_X1 FILLER_146_107 ();
 FILLCELL_X32 FILLER_146_128 ();
 FILLCELL_X8 FILLER_146_160 ();
 FILLCELL_X8 FILLER_146_188 ();
 FILLCELL_X1 FILLER_146_196 ();
 FILLCELL_X32 FILLER_146_202 ();
 FILLCELL_X32 FILLER_146_234 ();
 FILLCELL_X32 FILLER_146_266 ();
 FILLCELL_X16 FILLER_146_298 ();
 FILLCELL_X4 FILLER_146_314 ();
 FILLCELL_X1 FILLER_146_318 ();
 FILLCELL_X8 FILLER_146_337 ();
 FILLCELL_X1 FILLER_146_345 ();
 FILLCELL_X1 FILLER_146_394 ();
 FILLCELL_X8 FILLER_146_495 ();
 FILLCELL_X1 FILLER_146_503 ();
 FILLCELL_X16 FILLER_146_506 ();
 FILLCELL_X4 FILLER_146_522 ();
 FILLCELL_X2 FILLER_146_526 ();
 FILLCELL_X1 FILLER_146_553 ();
 FILLCELL_X2 FILLER_146_574 ();
 FILLCELL_X1 FILLER_146_586 ();
 FILLCELL_X4 FILLER_146_589 ();
 FILLCELL_X1 FILLER_146_593 ();
 FILLCELL_X1 FILLER_146_613 ();
 FILLCELL_X1 FILLER_146_617 ();
 FILLCELL_X2 FILLER_146_628 ();
 FILLCELL_X1 FILLER_146_630 ();
 FILLCELL_X1 FILLER_146_632 ();
 FILLCELL_X1 FILLER_146_688 ();
 FILLCELL_X1 FILLER_146_705 ();
 FILLCELL_X1 FILLER_146_710 ();
 FILLCELL_X1 FILLER_146_713 ();
 FILLCELL_X2 FILLER_146_732 ();
 FILLCELL_X1 FILLER_146_805 ();
 FILLCELL_X4 FILLER_146_810 ();
 FILLCELL_X2 FILLER_146_840 ();
 FILLCELL_X32 FILLER_146_887 ();
 FILLCELL_X32 FILLER_146_919 ();
 FILLCELL_X4 FILLER_146_951 ();
 FILLCELL_X2 FILLER_146_971 ();
 FILLCELL_X2 FILLER_146_983 ();
 FILLCELL_X8 FILLER_146_1007 ();
 FILLCELL_X2 FILLER_146_1015 ();
 FILLCELL_X1 FILLER_146_1017 ();
 FILLCELL_X2 FILLER_146_1044 ();
 FILLCELL_X1 FILLER_146_1053 ();
 FILLCELL_X1 FILLER_146_1065 ();
 FILLCELL_X1 FILLER_146_1078 ();
 FILLCELL_X1 FILLER_146_1087 ();
 FILLCELL_X32 FILLER_146_1091 ();
 FILLCELL_X16 FILLER_146_1123 ();
 FILLCELL_X8 FILLER_146_1139 ();
 FILLCELL_X1 FILLER_146_1147 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X2 FILLER_147_321 ();
 FILLCELL_X1 FILLER_147_323 ();
 FILLCELL_X1 FILLER_147_340 ();
 FILLCELL_X2 FILLER_147_343 ();
 FILLCELL_X1 FILLER_147_345 ();
 FILLCELL_X4 FILLER_147_348 ();
 FILLCELL_X4 FILLER_147_356 ();
 FILLCELL_X2 FILLER_147_360 ();
 FILLCELL_X1 FILLER_147_362 ();
 FILLCELL_X8 FILLER_147_365 ();
 FILLCELL_X2 FILLER_147_373 ();
 FILLCELL_X1 FILLER_147_375 ();
 FILLCELL_X8 FILLER_147_410 ();
 FILLCELL_X2 FILLER_147_418 ();
 FILLCELL_X4 FILLER_147_424 ();
 FILLCELL_X2 FILLER_147_476 ();
 FILLCELL_X1 FILLER_147_478 ();
 FILLCELL_X8 FILLER_147_481 ();
 FILLCELL_X4 FILLER_147_534 ();
 FILLCELL_X1 FILLER_147_538 ();
 FILLCELL_X4 FILLER_147_557 ();
 FILLCELL_X2 FILLER_147_561 ();
 FILLCELL_X1 FILLER_147_563 ();
 FILLCELL_X4 FILLER_147_584 ();
 FILLCELL_X2 FILLER_147_588 ();
 FILLCELL_X8 FILLER_147_592 ();
 FILLCELL_X1 FILLER_147_600 ();
 FILLCELL_X2 FILLER_147_603 ();
 FILLCELL_X1 FILLER_147_615 ();
 FILLCELL_X4 FILLER_147_636 ();
 FILLCELL_X2 FILLER_147_640 ();
 FILLCELL_X2 FILLER_147_646 ();
 FILLCELL_X1 FILLER_147_648 ();
 FILLCELL_X1 FILLER_147_655 ();
 FILLCELL_X2 FILLER_147_660 ();
 FILLCELL_X8 FILLER_147_680 ();
 FILLCELL_X1 FILLER_147_688 ();
 FILLCELL_X16 FILLER_147_693 ();
 FILLCELL_X1 FILLER_147_717 ();
 FILLCELL_X4 FILLER_147_726 ();
 FILLCELL_X1 FILLER_147_730 ();
 FILLCELL_X16 FILLER_147_733 ();
 FILLCELL_X8 FILLER_147_749 ();
 FILLCELL_X1 FILLER_147_757 ();
 FILLCELL_X4 FILLER_147_780 ();
 FILLCELL_X4 FILLER_147_794 ();
 FILLCELL_X1 FILLER_147_798 ();
 FILLCELL_X2 FILLER_147_852 ();
 FILLCELL_X32 FILLER_147_871 ();
 FILLCELL_X32 FILLER_147_903 ();
 FILLCELL_X16 FILLER_147_935 ();
 FILLCELL_X4 FILLER_147_951 ();
 FILLCELL_X4 FILLER_147_965 ();
 FILLCELL_X2 FILLER_147_969 ();
 FILLCELL_X1 FILLER_147_971 ();
 FILLCELL_X16 FILLER_147_976 ();
 FILLCELL_X32 FILLER_147_994 ();
 FILLCELL_X4 FILLER_147_1026 ();
 FILLCELL_X2 FILLER_147_1030 ();
 FILLCELL_X1 FILLER_147_1032 ();
 FILLCELL_X1 FILLER_147_1059 ();
 FILLCELL_X32 FILLER_147_1092 ();
 FILLCELL_X16 FILLER_147_1124 ();
 FILLCELL_X8 FILLER_147_1140 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X8 FILLER_148_321 ();
 FILLCELL_X4 FILLER_148_329 ();
 FILLCELL_X1 FILLER_148_333 ();
 FILLCELL_X1 FILLER_148_338 ();
 FILLCELL_X1 FILLER_148_355 ();
 FILLCELL_X4 FILLER_148_372 ();
 FILLCELL_X1 FILLER_148_380 ();
 FILLCELL_X1 FILLER_148_385 ();
 FILLCELL_X4 FILLER_148_397 ();
 FILLCELL_X1 FILLER_148_405 ();
 FILLCELL_X1 FILLER_148_410 ();
 FILLCELL_X1 FILLER_148_417 ();
 FILLCELL_X1 FILLER_148_434 ();
 FILLCELL_X1 FILLER_148_441 ();
 FILLCELL_X1 FILLER_148_444 ();
 FILLCELL_X1 FILLER_148_503 ();
 FILLCELL_X2 FILLER_148_520 ();
 FILLCELL_X2 FILLER_148_551 ();
 FILLCELL_X1 FILLER_148_553 ();
 FILLCELL_X8 FILLER_148_568 ();
 FILLCELL_X4 FILLER_148_576 ();
 FILLCELL_X4 FILLER_148_590 ();
 FILLCELL_X1 FILLER_148_594 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X2 FILLER_148_636 ();
 FILLCELL_X2 FILLER_148_642 ();
 FILLCELL_X4 FILLER_148_660 ();
 FILLCELL_X1 FILLER_148_664 ();
 FILLCELL_X2 FILLER_148_673 ();
 FILLCELL_X1 FILLER_148_675 ();
 FILLCELL_X1 FILLER_148_680 ();
 FILLCELL_X1 FILLER_148_683 ();
 FILLCELL_X2 FILLER_148_698 ();
 FILLCELL_X1 FILLER_148_702 ();
 FILLCELL_X2 FILLER_148_739 ();
 FILLCELL_X4 FILLER_148_761 ();
 FILLCELL_X2 FILLER_148_785 ();
 FILLCELL_X1 FILLER_148_787 ();
 FILLCELL_X4 FILLER_148_823 ();
 FILLCELL_X4 FILLER_148_870 ();
 FILLCELL_X2 FILLER_148_874 ();
 FILLCELL_X32 FILLER_148_903 ();
 FILLCELL_X32 FILLER_148_935 ();
 FILLCELL_X32 FILLER_148_967 ();
 FILLCELL_X32 FILLER_148_999 ();
 FILLCELL_X8 FILLER_148_1031 ();
 FILLCELL_X2 FILLER_148_1039 ();
 FILLCELL_X1 FILLER_148_1041 ();
 FILLCELL_X8 FILLER_148_1045 ();
 FILLCELL_X2 FILLER_148_1053 ();
 FILLCELL_X32 FILLER_148_1058 ();
 FILLCELL_X32 FILLER_148_1090 ();
 FILLCELL_X16 FILLER_148_1122 ();
 FILLCELL_X8 FILLER_148_1138 ();
 FILLCELL_X2 FILLER_148_1146 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X4 FILLER_149_321 ();
 FILLCELL_X2 FILLER_149_325 ();
 FILLCELL_X1 FILLER_149_327 ();
 FILLCELL_X1 FILLER_149_346 ();
 FILLCELL_X1 FILLER_149_369 ();
 FILLCELL_X1 FILLER_149_390 ();
 FILLCELL_X1 FILLER_149_410 ();
 FILLCELL_X4 FILLER_149_449 ();
 FILLCELL_X2 FILLER_149_453 ();
 FILLCELL_X8 FILLER_149_459 ();
 FILLCELL_X2 FILLER_149_467 ();
 FILLCELL_X2 FILLER_149_473 ();
 FILLCELL_X1 FILLER_149_475 ();
 FILLCELL_X2 FILLER_149_503 ();
 FILLCELL_X1 FILLER_149_505 ();
 FILLCELL_X1 FILLER_149_534 ();
 FILLCELL_X8 FILLER_149_537 ();
 FILLCELL_X8 FILLER_149_549 ();
 FILLCELL_X1 FILLER_149_557 ();
 FILLCELL_X1 FILLER_149_565 ();
 FILLCELL_X2 FILLER_149_596 ();
 FILLCELL_X1 FILLER_149_601 ();
 FILLCELL_X1 FILLER_149_604 ();
 FILLCELL_X2 FILLER_149_608 ();
 FILLCELL_X2 FILLER_149_650 ();
 FILLCELL_X4 FILLER_149_656 ();
 FILLCELL_X1 FILLER_149_667 ();
 FILLCELL_X4 FILLER_149_752 ();
 FILLCELL_X2 FILLER_149_756 ();
 FILLCELL_X2 FILLER_149_760 ();
 FILLCELL_X1 FILLER_149_762 ();
 FILLCELL_X1 FILLER_149_803 ();
 FILLCELL_X4 FILLER_149_855 ();
 FILLCELL_X1 FILLER_149_859 ();
 FILLCELL_X32 FILLER_149_882 ();
 FILLCELL_X32 FILLER_149_914 ();
 FILLCELL_X32 FILLER_149_946 ();
 FILLCELL_X32 FILLER_149_978 ();
 FILLCELL_X32 FILLER_149_1010 ();
 FILLCELL_X32 FILLER_149_1042 ();
 FILLCELL_X32 FILLER_149_1074 ();
 FILLCELL_X32 FILLER_149_1106 ();
 FILLCELL_X8 FILLER_149_1138 ();
 FILLCELL_X2 FILLER_149_1146 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X1 FILLER_150_321 ();
 FILLCELL_X2 FILLER_150_338 ();
 FILLCELL_X1 FILLER_150_340 ();
 FILLCELL_X2 FILLER_150_347 ();
 FILLCELL_X1 FILLER_150_349 ();
 FILLCELL_X2 FILLER_150_395 ();
 FILLCELL_X1 FILLER_150_401 ();
 FILLCELL_X1 FILLER_150_406 ();
 FILLCELL_X2 FILLER_150_409 ();
 FILLCELL_X4 FILLER_150_415 ();
 FILLCELL_X2 FILLER_150_419 ();
 FILLCELL_X1 FILLER_150_425 ();
 FILLCELL_X1 FILLER_150_430 ();
 FILLCELL_X1 FILLER_150_435 ();
 FILLCELL_X1 FILLER_150_452 ();
 FILLCELL_X4 FILLER_150_472 ();
 FILLCELL_X2 FILLER_150_510 ();
 FILLCELL_X4 FILLER_150_514 ();
 FILLCELL_X2 FILLER_150_538 ();
 FILLCELL_X1 FILLER_150_540 ();
 FILLCELL_X2 FILLER_150_621 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X2 FILLER_150_668 ();
 FILLCELL_X4 FILLER_150_674 ();
 FILLCELL_X1 FILLER_150_678 ();
 FILLCELL_X4 FILLER_150_683 ();
 FILLCELL_X4 FILLER_150_691 ();
 FILLCELL_X1 FILLER_150_695 ();
 FILLCELL_X1 FILLER_150_712 ();
 FILLCELL_X1 FILLER_150_717 ();
 FILLCELL_X4 FILLER_150_722 ();
 FILLCELL_X2 FILLER_150_726 ();
 FILLCELL_X1 FILLER_150_728 ();
 FILLCELL_X8 FILLER_150_731 ();
 FILLCELL_X2 FILLER_150_739 ();
 FILLCELL_X2 FILLER_150_807 ();
 FILLCELL_X2 FILLER_150_821 ();
 FILLCELL_X1 FILLER_150_841 ();
 FILLCELL_X8 FILLER_150_846 ();
 FILLCELL_X1 FILLER_150_854 ();
 FILLCELL_X32 FILLER_150_877 ();
 FILLCELL_X32 FILLER_150_909 ();
 FILLCELL_X32 FILLER_150_941 ();
 FILLCELL_X32 FILLER_150_973 ();
 FILLCELL_X32 FILLER_150_1005 ();
 FILLCELL_X32 FILLER_150_1037 ();
 FILLCELL_X32 FILLER_150_1069 ();
 FILLCELL_X32 FILLER_150_1101 ();
 FILLCELL_X8 FILLER_150_1133 ();
 FILLCELL_X4 FILLER_150_1141 ();
 FILLCELL_X2 FILLER_150_1145 ();
 FILLCELL_X1 FILLER_150_1147 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X4 FILLER_151_321 ();
 FILLCELL_X1 FILLER_151_325 ();
 FILLCELL_X8 FILLER_151_328 ();
 FILLCELL_X2 FILLER_151_336 ();
 FILLCELL_X1 FILLER_151_373 ();
 FILLCELL_X1 FILLER_151_420 ();
 FILLCELL_X1 FILLER_151_439 ();
 FILLCELL_X2 FILLER_151_442 ();
 FILLCELL_X1 FILLER_151_458 ();
 FILLCELL_X8 FILLER_151_493 ();
 FILLCELL_X4 FILLER_151_501 ();
 FILLCELL_X2 FILLER_151_505 ();
 FILLCELL_X1 FILLER_151_507 ();
 FILLCELL_X1 FILLER_151_526 ();
 FILLCELL_X2 FILLER_151_581 ();
 FILLCELL_X8 FILLER_151_593 ();
 FILLCELL_X1 FILLER_151_601 ();
 FILLCELL_X1 FILLER_151_647 ();
 FILLCELL_X1 FILLER_151_653 ();
 FILLCELL_X1 FILLER_151_728 ();
 FILLCELL_X8 FILLER_151_733 ();
 FILLCELL_X4 FILLER_151_741 ();
 FILLCELL_X1 FILLER_151_745 ();
 FILLCELL_X32 FILLER_151_879 ();
 FILLCELL_X32 FILLER_151_911 ();
 FILLCELL_X32 FILLER_151_943 ();
 FILLCELL_X32 FILLER_151_975 ();
 FILLCELL_X32 FILLER_151_1007 ();
 FILLCELL_X32 FILLER_151_1039 ();
 FILLCELL_X32 FILLER_151_1071 ();
 FILLCELL_X32 FILLER_151_1103 ();
 FILLCELL_X8 FILLER_151_1135 ();
 FILLCELL_X4 FILLER_151_1143 ();
 FILLCELL_X1 FILLER_151_1147 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X8 FILLER_152_337 ();
 FILLCELL_X2 FILLER_152_345 ();
 FILLCELL_X2 FILLER_152_349 ();
 FILLCELL_X1 FILLER_152_355 ();
 FILLCELL_X1 FILLER_152_364 ();
 FILLCELL_X4 FILLER_152_373 ();
 FILLCELL_X8 FILLER_152_389 ();
 FILLCELL_X1 FILLER_152_397 ();
 FILLCELL_X1 FILLER_152_406 ();
 FILLCELL_X1 FILLER_152_427 ();
 FILLCELL_X2 FILLER_152_446 ();
 FILLCELL_X1 FILLER_152_448 ();
 FILLCELL_X1 FILLER_152_455 ();
 FILLCELL_X1 FILLER_152_460 ();
 FILLCELL_X4 FILLER_152_463 ();
 FILLCELL_X2 FILLER_152_469 ();
 FILLCELL_X2 FILLER_152_473 ();
 FILLCELL_X2 FILLER_152_479 ();
 FILLCELL_X1 FILLER_152_481 ();
 FILLCELL_X4 FILLER_152_486 ();
 FILLCELL_X1 FILLER_152_490 ();
 FILLCELL_X4 FILLER_152_495 ();
 FILLCELL_X4 FILLER_152_501 ();
 FILLCELL_X2 FILLER_152_505 ();
 FILLCELL_X4 FILLER_152_526 ();
 FILLCELL_X2 FILLER_152_547 ();
 FILLCELL_X1 FILLER_152_549 ();
 FILLCELL_X1 FILLER_152_555 ();
 FILLCELL_X1 FILLER_152_560 ();
 FILLCELL_X1 FILLER_152_565 ();
 FILLCELL_X2 FILLER_152_628 ();
 FILLCELL_X1 FILLER_152_630 ();
 FILLCELL_X1 FILLER_152_632 ();
 FILLCELL_X1 FILLER_152_636 ();
 FILLCELL_X4 FILLER_152_644 ();
 FILLCELL_X1 FILLER_152_652 ();
 FILLCELL_X1 FILLER_152_677 ();
 FILLCELL_X1 FILLER_152_680 ();
 FILLCELL_X2 FILLER_152_709 ();
 FILLCELL_X8 FILLER_152_713 ();
 FILLCELL_X2 FILLER_152_721 ();
 FILLCELL_X4 FILLER_152_739 ();
 FILLCELL_X2 FILLER_152_743 ();
 FILLCELL_X2 FILLER_152_796 ();
 FILLCELL_X1 FILLER_152_798 ();
 FILLCELL_X2 FILLER_152_814 ();
 FILLCELL_X1 FILLER_152_816 ();
 FILLCELL_X1 FILLER_152_828 ();
 FILLCELL_X2 FILLER_152_840 ();
 FILLCELL_X1 FILLER_152_842 ();
 FILLCELL_X2 FILLER_152_846 ();
 FILLCELL_X2 FILLER_152_851 ();
 FILLCELL_X32 FILLER_152_873 ();
 FILLCELL_X32 FILLER_152_905 ();
 FILLCELL_X32 FILLER_152_937 ();
 FILLCELL_X32 FILLER_152_969 ();
 FILLCELL_X32 FILLER_152_1001 ();
 FILLCELL_X32 FILLER_152_1033 ();
 FILLCELL_X32 FILLER_152_1065 ();
 FILLCELL_X32 FILLER_152_1097 ();
 FILLCELL_X16 FILLER_152_1129 ();
 FILLCELL_X2 FILLER_152_1145 ();
 FILLCELL_X1 FILLER_152_1147 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X4 FILLER_153_321 ();
 FILLCELL_X8 FILLER_153_327 ();
 FILLCELL_X4 FILLER_153_335 ();
 FILLCELL_X2 FILLER_153_339 ();
 FILLCELL_X2 FILLER_153_357 ();
 FILLCELL_X1 FILLER_153_359 ();
 FILLCELL_X1 FILLER_153_414 ();
 FILLCELL_X1 FILLER_153_417 ();
 FILLCELL_X2 FILLER_153_448 ();
 FILLCELL_X1 FILLER_153_450 ();
 FILLCELL_X2 FILLER_153_519 ();
 FILLCELL_X4 FILLER_153_607 ();
 FILLCELL_X4 FILLER_153_694 ();
 FILLCELL_X2 FILLER_153_717 ();
 FILLCELL_X2 FILLER_153_751 ();
 FILLCELL_X1 FILLER_153_755 ();
 FILLCELL_X1 FILLER_153_762 ();
 FILLCELL_X2 FILLER_153_765 ();
 FILLCELL_X1 FILLER_153_772 ();
 FILLCELL_X2 FILLER_153_804 ();
 FILLCELL_X1 FILLER_153_806 ();
 FILLCELL_X1 FILLER_153_832 ();
 FILLCELL_X1 FILLER_153_859 ();
 FILLCELL_X32 FILLER_153_882 ();
 FILLCELL_X32 FILLER_153_914 ();
 FILLCELL_X32 FILLER_153_946 ();
 FILLCELL_X32 FILLER_153_978 ();
 FILLCELL_X32 FILLER_153_1010 ();
 FILLCELL_X32 FILLER_153_1042 ();
 FILLCELL_X32 FILLER_153_1074 ();
 FILLCELL_X32 FILLER_153_1106 ();
 FILLCELL_X8 FILLER_153_1138 ();
 FILLCELL_X2 FILLER_153_1146 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X16 FILLER_154_97 ();
 FILLCELL_X8 FILLER_154_113 ();
 FILLCELL_X2 FILLER_154_121 ();
 FILLCELL_X32 FILLER_154_130 ();
 FILLCELL_X32 FILLER_154_162 ();
 FILLCELL_X32 FILLER_154_194 ();
 FILLCELL_X32 FILLER_154_226 ();
 FILLCELL_X32 FILLER_154_258 ();
 FILLCELL_X32 FILLER_154_290 ();
 FILLCELL_X8 FILLER_154_322 ();
 FILLCELL_X2 FILLER_154_332 ();
 FILLCELL_X4 FILLER_154_354 ();
 FILLCELL_X2 FILLER_154_358 ();
 FILLCELL_X8 FILLER_154_364 ();
 FILLCELL_X2 FILLER_154_372 ();
 FILLCELL_X1 FILLER_154_376 ();
 FILLCELL_X4 FILLER_154_385 ();
 FILLCELL_X4 FILLER_154_403 ();
 FILLCELL_X1 FILLER_154_407 ();
 FILLCELL_X2 FILLER_154_421 ();
 FILLCELL_X2 FILLER_154_440 ();
 FILLCELL_X2 FILLER_154_446 ();
 FILLCELL_X1 FILLER_154_454 ();
 FILLCELL_X2 FILLER_154_469 ();
 FILLCELL_X4 FILLER_154_483 ();
 FILLCELL_X1 FILLER_154_491 ();
 FILLCELL_X2 FILLER_154_496 ();
 FILLCELL_X2 FILLER_154_502 ();
 FILLCELL_X2 FILLER_154_509 ();
 FILLCELL_X1 FILLER_154_511 ();
 FILLCELL_X1 FILLER_154_516 ();
 FILLCELL_X4 FILLER_154_541 ();
 FILLCELL_X4 FILLER_154_555 ();
 FILLCELL_X4 FILLER_154_562 ();
 FILLCELL_X2 FILLER_154_589 ();
 FILLCELL_X2 FILLER_154_599 ();
 FILLCELL_X1 FILLER_154_607 ();
 FILLCELL_X1 FILLER_154_611 ();
 FILLCELL_X1 FILLER_154_635 ();
 FILLCELL_X1 FILLER_154_668 ();
 FILLCELL_X1 FILLER_154_673 ();
 FILLCELL_X2 FILLER_154_678 ();
 FILLCELL_X2 FILLER_154_683 ();
 FILLCELL_X2 FILLER_154_688 ();
 FILLCELL_X1 FILLER_154_690 ();
 FILLCELL_X4 FILLER_154_707 ();
 FILLCELL_X1 FILLER_154_711 ();
 FILLCELL_X2 FILLER_154_775 ();
 FILLCELL_X1 FILLER_154_855 ();
 FILLCELL_X32 FILLER_154_890 ();
 FILLCELL_X32 FILLER_154_922 ();
 FILLCELL_X32 FILLER_154_954 ();
 FILLCELL_X32 FILLER_154_986 ();
 FILLCELL_X32 FILLER_154_1018 ();
 FILLCELL_X32 FILLER_154_1050 ();
 FILLCELL_X32 FILLER_154_1082 ();
 FILLCELL_X32 FILLER_154_1114 ();
 FILLCELL_X2 FILLER_154_1146 ();
endmodule
