module dadda11(a, b, t1, t2);
output wire [21:0] t1, t2;
input wire [10:0] a, b;
wire wire_1, wire_2;
wire wire_3, wire_4;
wire wire_5, wire_6;
wire wire_7, wire_8;
wire wire_9, wire_10;
wire wire_11, wire_12;
wire wire_13, wire_14;
wire wire_15, wire_16;
wire wire_17, wire_18;
wire wire_19, wire_20;
wire wire_21, wire_22;
wire wire_23, wire_24;
wire wire_25, wire_26;
wire wire_27, wire_28;
wire wire_29, wire_30;
wire wire_31, wire_32;
wire wire_33, wire_34;
wire wire_35, wire_36;
wire wire_37, wire_38;
wire wire_39, wire_40;
wire wire_41, wire_42;
wire wire_43, wire_44;
wire wire_45, wire_46;
wire wire_47, wire_48;
wire wire_49, wire_50;
wire wire_51, wire_52;
wire wire_53, wire_54;
wire wire_55, wire_56;
wire wire_57, wire_58;
wire wire_59, wire_60;
wire wire_61, wire_62;
wire wire_63, wire_64;
wire wire_65, wire_66;
wire wire_67, wire_68;
wire wire_69, wire_70;
wire wire_71, wire_72;
wire wire_73, wire_74;
wire wire_75, wire_76;
wire wire_77, wire_78;
wire wire_79, wire_80;
wire wire_81, wire_82;
wire wire_83, wire_84;
wire wire_85, wire_86;
wire wire_87, wire_88;
wire wire_89, wire_90;
wire wire_91, wire_92;
wire wire_93, wire_94;
wire wire_95, wire_96;
wire wire_97, wire_98;
wire wire_99, wire_100;
wire wire_101, wire_102;
wire wire_103, wire_104;
wire wire_105, wire_106;
wire wire_107, wire_108;
wire wire_109, wire_110;
wire wire_111, wire_112;
wire wire_113, wire_114;
wire wire_115, wire_116;
wire wire_117, wire_118;
wire wire_119, wire_120;
wire wire_121, wire_122;
wire wire_123, wire_124;
wire wire_125, wire_126;
wire wire_127, wire_128;
wire wire_129, wire_130;
wire wire_131, wire_132;
wire wire_133, wire_134;
wire wire_135, wire_136;
wire wire_137, wire_138;
wire wire_139, wire_140;
wire wire_141, wire_142;
wire wire_143, wire_144;
wire wire_145, wire_146;
wire wire_147, wire_148;
wire wire_149, wire_150;
wire wire_151, wire_152;
wire wire_153, wire_154;
wire wire_155, wire_156;
wire wire_157, wire_158;
wire wire_159, wire_160;
wire wire_161, wire_162;
wire wire_163, wire_164;
wire wire_165, wire_166;
wire wire_167, wire_168;
wire wire_169, wire_170;
wire wire_171, wire_172;
wire wire_173, wire_174;
wire wire_175, wire_176;
wire wire_177, wire_178;
wire wire_179, wire_180;
assign {{ wire_1, wire_2 }} = (a[0] & b[9]) + (a[1] & b[8]);
assign {{ wire_3, wire_4 }} = (a[0] & b[10]) + (a[1] & b[9]) + (a[2] & b[8]);
assign {{ wire_5, wire_6 }} = (a[3] & b[7]) + (a[4] & b[6]);
assign {{ wire_7, wire_8 }} = (a[1] & b[10]) + (a[2] & b[9]) + (a[3] & b[8]);
assign {{ wire_9, wire_10 }} = (a[4] & b[7]) + (a[5] & b[6]);
assign {{ wire_11, wire_12 }} = (a[2] & b[10]) + (a[3] & b[9]) + (a[4] & b[8]);
assign {{ wire_13, wire_14 }} = (a[0] & b[6]) + (a[1] & b[5]);
assign {{ wire_15, wire_16 }} = (a[0] & b[7]) + (a[1] & b[6]) + (a[2] & b[5]);
assign {{ wire_17, wire_18 }} = (a[3] & b[4]) + (a[4] & b[3]);
assign {{ wire_19, wire_20 }} = (a[0] & b[8]) + (a[1] & b[7]) + (a[2] & b[6]);
assign {{ wire_21, wire_22 }} = (a[3] & b[5]) + (a[4] & b[4]) + (a[5] & b[3]);
assign {{ wire_23, wire_24 }} = (a[6] & b[2]) + (a[7] & b[1]);
assign {{ wire_25, wire_26 }} = (a[2] & b[7]) + (a[3] & b[6]) + (a[4] & b[5]);
assign {{ wire_27, wire_28 }} = (a[5] & b[4]) + (a[6] & b[3]) + (a[7] & b[2]);
assign {{ wire_29, wire_30 }} = (a[8] & b[1]) + (a[9] & b[0]) + wire_2;
assign {{ wire_31, wire_32 }} = (a[5] & b[5]) + (a[6] & b[4]) + (a[7] & b[3]);
assign {{ wire_33, wire_34 }} = (a[8] & b[2]) + (a[9] & b[1]) + (a[10] & b[0]);
assign {{ wire_35, wire_36 }} = wire_1 + wire_4 + wire_6;
assign {{ wire_37, wire_38 }} = (a[6] & b[5]) + (a[7] & b[4]) + (a[8] & b[3]);
assign {{ wire_39, wire_40 }} = (a[9] & b[2]) + (a[10] & b[1]) + wire_3;
assign {{ wire_41, wire_42 }} = wire_5 + wire_8 + wire_10;
assign {{ wire_43, wire_44 }} = (a[5] & b[7]) + (a[6] & b[6]) + (a[7] & b[5]);
assign {{ wire_45, wire_46 }} = (a[8] & b[4]) + (a[9] & b[3]) + (a[10] & b[2]);
assign {{ wire_47, wire_48 }} = wire_7 + wire_9 + wire_12;
assign {{ wire_49, wire_50 }} = (a[3] & b[10]) + (a[4] & b[9]) + (a[5] & b[8]);
assign {{ wire_51, wire_52 }} = (a[6] & b[7]) + (a[7] & b[6]) + (a[8] & b[5]);
assign {{ wire_53, wire_54 }} = (a[9] & b[4]) + (a[10] & b[3]) + wire_11;
assign {{ wire_55, wire_56 }} = (a[4] & b[10]) + (a[5] & b[9]) + (a[6] & b[8]);
assign {{ wire_57, wire_58 }} = (a[7] & b[7]) + (a[8] & b[6]) + (a[9] & b[5]);
assign {{ wire_59, wire_60 }} = (a[5] & b[10]) + (a[6] & b[9]) + (a[7] & b[8]);
assign {{ wire_61, wire_62 }} = (a[0] & b[4]) + (a[1] & b[3]);
assign {{ wire_63, wire_64 }} = (a[0] & b[5]) + (a[1] & b[4]) + (a[2] & b[3]);
assign {{ wire_65, wire_66 }} = (a[3] & b[2]) + (a[4] & b[1]);
assign {{ wire_67, wire_68 }} = (a[2] & b[4]) + (a[3] & b[3]) + (a[4] & b[2]);
assign {{ wire_69, wire_70 }} = (a[5] & b[1]) + (a[6] & b[0]) + wire_14;
assign {{ wire_71, wire_72 }} = (a[5] & b[2]) + (a[6] & b[1]) + (a[7] & b[0]);
assign {{ wire_73, wire_74 }} = wire_13 + wire_16 + wire_18;
assign {{ wire_75, wire_76 }} = (a[8] & b[0]) + wire_15 + wire_17;
assign {{ wire_77, wire_78 }} = wire_20 + wire_22 + wire_24;
assign {{ wire_79, wire_80 }} = wire_19 + wire_21 + wire_23;
assign {{ wire_81, wire_82 }} = wire_26 + wire_28 + wire_30;
assign {{ wire_83, wire_84 }} = wire_25 + wire_27 + wire_29;
assign {{ wire_85, wire_86 }} = wire_32 + wire_34 + wire_36;
assign {{ wire_87, wire_88 }} = wire_31 + wire_33 + wire_35;
assign {{ wire_89, wire_90 }} = wire_38 + wire_40 + wire_42;
assign {{ wire_91, wire_92 }} = wire_37 + wire_39 + wire_41;
assign {{ wire_93, wire_94 }} = wire_44 + wire_46 + wire_48;
assign {{ wire_95, wire_96 }} = wire_43 + wire_45 + wire_47;
assign {{ wire_97, wire_98 }} = wire_50 + wire_52 + wire_54;
assign {{ wire_99, wire_100 }} = (a[10] & b[4]) + wire_49 + wire_51;
assign {{ wire_101, wire_102 }} = wire_53 + wire_56 + wire_58;
assign {{ wire_103, wire_104 }} = (a[8] & b[7]) + (a[9] & b[6]) + (a[10] & b[5]);
assign {{ wire_105, wire_106 }} = wire_55 + wire_57 + wire_60;
assign {{ wire_107, wire_108 }} = (a[6] & b[10]) + (a[7] & b[9]) + (a[8] & b[8]);
assign {{ wire_109, wire_110 }} = (a[9] & b[7]) + (a[10] & b[6]) + wire_59;
assign {{ wire_111, wire_112 }} = (a[7] & b[10]) + (a[8] & b[9]) + (a[9] & b[8]);
assign {{ wire_113, wire_114 }} = (a[0] & b[3]) + (a[1] & b[2]);
assign {{ wire_115, wire_116 }} = (a[2] & b[2]) + (a[3] & b[1]) + (a[4] & b[0]);
assign {{ wire_117, wire_118 }} = (a[5] & b[0]) + wire_61 + wire_64;
assign {{ wire_119, wire_120 }} = wire_63 + wire_65 + wire_68;
assign {{ wire_121, wire_122 }} = wire_67 + wire_69 + wire_72;
assign {{ wire_123, wire_124 }} = wire_71 + wire_73 + wire_76;
assign {{ wire_125, wire_126 }} = wire_75 + wire_77 + wire_80;
assign {{ wire_127, wire_128 }} = wire_79 + wire_81 + wire_84;
assign {{ wire_129, wire_130 }} = wire_83 + wire_85 + wire_88;
assign {{ wire_131, wire_132 }} = wire_87 + wire_89 + wire_92;
assign {{ wire_133, wire_134 }} = wire_91 + wire_93 + wire_96;
assign {{ wire_135, wire_136 }} = wire_95 + wire_97 + wire_100;
assign {{ wire_137, wire_138 }} = wire_99 + wire_101 + wire_104;
assign {{ wire_139, wire_140 }} = wire_103 + wire_105 + wire_108;
assign {{ wire_141, wire_142 }} = (a[10] & b[7]) + wire_107 + wire_109;
assign {{ wire_143, wire_144 }} = (a[8] & b[10]) + (a[9] & b[9]) + (a[10] & b[8]);
assign {{ wire_145, wire_146 }} = (a[0] & b[2]) + (a[1] & b[1]);
assign {{ wire_147, wire_148 }} = (a[2] & b[1]) + (a[3] & b[0]) + wire_114;
assign {{ wire_149, wire_150 }} = wire_62 + wire_113 + wire_116;
assign {{ wire_151, wire_152 }} = wire_66 + wire_115 + wire_118;
assign {{ wire_153, wire_154 }} = wire_70 + wire_117 + wire_120;
assign {{ wire_155, wire_156 }} = wire_74 + wire_119 + wire_122;
assign {{ wire_157, wire_158 }} = wire_78 + wire_121 + wire_124;
assign {{ wire_159, wire_160 }} = wire_82 + wire_123 + wire_126;
assign {{ wire_161, wire_162 }} = wire_86 + wire_125 + wire_128;
assign {{ wire_163, wire_164 }} = wire_90 + wire_127 + wire_130;
assign {{ wire_165, wire_166 }} = wire_94 + wire_129 + wire_132;
assign {{ wire_167, wire_168 }} = wire_98 + wire_131 + wire_134;
assign {{ wire_169, wire_170 }} = wire_102 + wire_133 + wire_136;
assign {{ wire_171, wire_172 }} = wire_106 + wire_135 + wire_138;
assign {{ wire_173, wire_174 }} = wire_110 + wire_137 + wire_140;
assign {{ wire_175, wire_176 }} = wire_112 + wire_139 + wire_142;
assign {{ wire_177, wire_178 }} = wire_111 + wire_141 + wire_144;
assign {{ wire_179, wire_180 }} = (a[9] & b[10]) + (a[10] & b[9]) + wire_143;
assign t1 = {(a[10] & b[10]),wire_177,wire_175,wire_173,wire_171,wire_169,wire_167,wire_165,wire_163,wire_161,wire_159,wire_157,wire_155,wire_153,wire_151,wire_149,wire_147,wire_145,(a[2] & b[0]),(a[0] & b[1]),(a[0] & b[0])};
assign t2 = {wire_179,wire_180,wire_178,wire_176,wire_174,wire_172,wire_170,wire_168,wire_166,wire_164,wire_162,wire_160,wire_158,wire_156,wire_154,wire_152,wire_150,wire_148,wire_146,(a[1] & b[0]),1'b0};
endmodule
